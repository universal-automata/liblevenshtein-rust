(** * Acceptance Criteria for Levenshtein Automata

    This module defines when a state is accepting and when the automaton
    accepts a dictionary word.

    Part of: Liblevenshtein.Core.Automaton

    Rust Reference: src/transducer/state.rs

    Key Definitions:
    - is_final: Whether an automaton state is final (accepting)
    - automaton_run: Run automaton on a dictionary word
    - automaton_accepts: Whether automaton accepts a dictionary word
    - accepting_distance: Minimum edit distance for accepted words

    Key Theorems:
    - final_state_characterization
    - accepting_distance_correct
    - run_deterministic
*)

From Stdlib Require Import Arith Bool List Nat Lia.
Import ListNotations.

From Liblevenshtein.Core Require Import Core.Definitions.
From Liblevenshtein.Core Require Import Automaton.Position.
From Liblevenshtein.Core Require Import Automaton.State.
From Liblevenshtein.Core Require Import Automaton.Transition.

(** * Final State Predicate *)

(** A position is final if it has consumed all of the query
    (term_index >= query_length). The remaining query characters
    are deletions, contributing to the error count. *)
Definition position_is_final (qlen : nat) (p : Position) : bool :=
  qlen <=? term_index p.

(** A state is final if it contains at least one final position.
    The minimum error count among final positions gives the edit distance. *)
Definition state_is_final (s : State) : bool :=
  existsb (position_is_final (query_length s)) (positions s).

(** * Accepting Distance *)

(** For a final position at term_index i (where i >= qlen),
    the total edit distance includes the position's errors plus
    any remaining deletions (i - qlen). But actually for our encoding,
    the num_errors already accounts for the path taken, so we just
    need to ensure the position can reach the end of the query. *)

(** Get the minimum error count among final positions *)
Definition final_position_distance (qlen : nat) (p : Position) : option nat :=
  if position_is_final qlen p then
    (* Distance = errors + remaining query chars to delete *)
    Some (num_errors p)
  else
    None.

Fixpoint min_option (a b : option nat) : option nat :=
  match a, b with
  | None, None => None
  | Some x, None => Some x
  | None, Some y => Some y
  | Some x, Some y => Some (min x y)
  end.

Definition state_accepting_distance (s : State) : option nat :=
  fold_right (fun p acc =>
    min_option (final_position_distance (query_length s) p) acc
  ) None (positions s).

(** * Automaton Run *)

(** Run the automaton on a dictionary word, returning the final state (or None if dead) *)
Fixpoint automaton_run (alg : Algorithm) (query : list Char) (n : nat)
                       (dict : list Char) (s : State) : option State :=
  match dict with
  | [] => Some s  (* End of dictionary word, return current state *)
  | c :: rest =>
      match transition_state alg s c query n with
      | None => None  (* Dead state *)
      | Some s' => automaton_run alg query n rest s'
      end
  end.

(** Run from initial state *)
Definition automaton_run_from_initial (alg : Algorithm) (query : list Char)
                                       (n : nat) (dict : list Char) : option State :=
  let qlen := length query in
  let init := initial_state alg qlen in
  (* First apply epsilon closure to initial state for delete operations *)
  let init_closed :=
    mkState (epsilon_closure (positions init) n qlen) alg qlen in
  automaton_run alg query n dict init_closed.

(** * Acceptance *)

(** Automaton accepts a dictionary word if the final state is accepting *)
Definition automaton_accepts (alg : Algorithm) (query : list Char)
                              (n : nat) (dict : list Char) : bool :=
  match automaton_run_from_initial alg query n dict with
  | None => false
  | Some final_state => state_is_final final_state
  end.

(** Get the accepting distance if the automaton accepts *)
Definition automaton_distance (alg : Algorithm) (query : list Char)
                               (n : nat) (dict : list Char) : option nat :=
  match automaton_run_from_initial alg query n dict with
  | None => None
  | Some final_state => state_accepting_distance final_state
  end.

(** * Properties *)

(** Final position characterization *)
Lemma position_final_iff : forall qlen p,
  position_is_final qlen p = true <-> qlen <= term_index p.
Proof.
  intros qlen p.
  unfold position_is_final.
  rewrite Nat.leb_le.
  reflexivity.
Qed.

(** State finality implies contains final position *)
Lemma state_final_has_final_position : forall s,
  state_is_final s = true ->
  exists p, In p (positions s) /\ position_is_final (query_length s) p = true.
Proof.
  intros s Hfinal.
  unfold state_is_final in Hfinal.
  rewrite existsb_exists in Hfinal.
  exact Hfinal.
Qed.

(** Helper: fold_right with min_option returns Some means some element was Some *)
Lemma fold_min_option_some_aux : forall {A} (f : A -> option nat) (l : list A) d,
  fold_right (fun x acc => min_option (f x) acc) None l = Some d ->
  exists a, In a l /\ exists d', f a = Some d' /\ d' >= d.
Proof.
  intros A f l. revert f.
  induction l as [| x xs IH]; intros f d Hfold.
  - simpl in Hfold. discriminate.
  - simpl in Hfold.
    set (rest := fold_right (fun x acc => min_option (f x) acc) None xs) in *.
    destruct (f x) as [dx|] eqn:Hfx; destruct rest as [dxs|] eqn:Hrest.
    + (* f x = Some dx, rest = Some dxs *)
      simpl in Hfold.
      assert (Hd : d = min dx dxs) by (inversion Hfold; reflexivity).
      destruct (Nat.min_dec dx dxs) as [Hmin | Hmin].
      * (* dx is min *)
        exists x. split; [left; reflexivity |].
        exists dx. split; [exact Hfx |].
        subst. rewrite Hmin. lia.
      * (* dxs is min *)
        unfold rest in Hrest.
        specialize (IH f dxs Hrest).
        destruct IH as [a [Hin [d' [Hfa Hge]]]].
        exists a. split; [right; exact Hin |].
        exists d'. split; [exact Hfa |].
        subst. rewrite Hmin. lia.
    + (* f x = Some dx, rest = None *)
      simpl in Hfold.
      assert (Hd : d = dx) by (inversion Hfold; reflexivity). subst.
      exists x. split; [left; reflexivity |].
      exists dx. split; [exact Hfx | lia].
    + (* f x = None, rest = Some dxs *)
      simpl in Hfold.
      assert (Hd : d = dxs) by (inversion Hfold; reflexivity). subst.
      unfold rest in Hrest.
      specialize (IH f dxs Hrest).
      destruct IH as [a [Hin [d' [Hfa Hge]]]].
      exists a. split; [right; exact Hin |].
      exists d'. split; [exact Hfa | exact Hge].
    + (* f x = None, rest = None *)
      simpl in Hfold. discriminate.
Qed.

Lemma fold_min_option_some : forall {A} (f : A -> option nat) (l : list A) d,
  fold_right (fun x acc => min_option (f x) acc) None l = Some d ->
  exists a, In a l /\ exists d', f a = Some d' /\ d' >= d.
Proof.
  intros A. exact (fold_min_option_some_aux (A := A)).
Qed.

(** The minimum is exactly achieved by some element *)
Lemma fold_min_option_achieves : forall {A} (f : A -> option nat) (l : list A) d,
  fold_right (fun x acc => min_option (f x) acc) None l = Some d ->
  exists a, In a l /\ f a = Some d.
Proof.
  intros A f l. revert f.
  induction l as [| x xs IH]; intros f d Hfold.
  - simpl in Hfold. discriminate.
  - simpl in Hfold.
    set (rest := fold_right (fun x acc => min_option (f x) acc) None xs) in *.
    destruct (f x) as [dx|] eqn:Hfx; destruct rest as [dr|] eqn:Hrest.
    + (* f x = Some dx, rest = Some dr *)
      simpl in Hfold.
      assert (Hd : d = min dx dr) by (inversion Hfold; reflexivity).
      destruct (Nat.min_dec dx dr) as [Hmin | Hmin].
      * (* dx <= dr, so d = dx *)
        subst d. rewrite Hmin.
        exists x. split; [left; reflexivity | exact Hfx].
      * (* dr < dx, so d = dr *)
        subst d. rewrite Hmin.
        unfold rest in Hrest.
        specialize (IH f dr Hrest).
        destruct IH as [a [Hin Ha]].
        exists a. split; [right; exact Hin | exact Ha].
    + (* f x = Some dx, rest = None *)
      simpl in Hfold.
      assert (Hd : d = dx) by (inversion Hfold; reflexivity). subst d.
      exists x. split; [left; reflexivity | exact Hfx].
    + (* f x = None, rest = Some dr *)
      simpl in Hfold.
      assert (Hd : d = dr) by (inversion Hfold; reflexivity). subst d.
      unfold rest in Hrest.
      specialize (IH f dr Hrest).
      destruct IH as [a [Hin Ha]].
      exists a. split; [right; exact Hin | exact Ha].
    + (* f x = None, rest = None *)
      simpl in Hfold. discriminate.
Qed.

(** Accepting distance is exactly achieved by some final position *)
Lemma accepting_distance_achieves : forall s d,
  state_accepting_distance s = Some d ->
  exists p, In p (positions s) /\
            position_is_final (query_length s) p = true /\
            num_errors p = d.
Proof.
  intros s d Hdist.
  unfold state_accepting_distance in Hdist.
  apply fold_min_option_achieves in Hdist.
  destruct Hdist as [p [Hin Hfpd]].
  unfold final_position_distance in Hfpd.
  destruct (position_is_final (query_length s) p) eqn:Hfinal.
  - inversion Hfpd.
    exists p. split; [exact Hin |]. split; [exact Hfinal | reflexivity].
  - discriminate.
Qed.

(** Accepting distance is achieved by some final position *)
Lemma accepting_distance_is_min : forall s d,
  state_accepting_distance s = Some d ->
  exists p, In p (positions s) /\
            position_is_final (query_length s) p = true /\
            num_errors p >= d.
Proof.
  intros s d Hdist.
  unfold state_accepting_distance in Hdist.
  apply fold_min_option_some in Hdist.
  destruct Hdist as [p [Hin [d' [Hfpd Hge]]]].
  unfold final_position_distance in Hfpd.
  destruct (position_is_final (query_length s) p) eqn:Hfinal.
  - inversion Hfpd. subst.
    exists p. split; [exact Hin |]. split; [exact Hfinal | exact Hge].
  - discriminate.
Qed.

(** Run is deterministic *)
Lemma run_deterministic : forall alg query n dict s s1 s2,
  automaton_run alg query n dict s = Some s1 ->
  automaton_run alg query n dict s = Some s2 ->
  s1 = s2.
Proof.
  intros alg query n dict s s1 s2 H1 H2.
  rewrite H1 in H2.
  inversion H2.
  reflexivity.
Qed.

(** Empty dictionary word: final state is initial state *)
Lemma run_empty_dict : forall alg query n s,
  automaton_run alg query n [] s = Some s.
Proof.
  intros alg query n s.
  simpl. reflexivity.
Qed.

(** * Helper Lemmas for Distance *)

(** If a position has term_index = qlen and e errors, distance is e *)
Lemma final_position_at_qlen : forall qlen i e s,
  i = qlen ->
  position_is_final qlen (mkPosition i e s) = true.
Proof.
  intros qlen i e s Heq.
  subst. unfold position_is_final. simpl.
  rewrite Nat.leb_refl. reflexivity.
Qed.

(** If a position has term_index > qlen, it's also final *)
Lemma final_position_past_qlen : forall qlen i e s,
  i > qlen ->
  position_is_final qlen (mkPosition i e s) = true.
Proof.
  intros qlen i e s Hgt.
  unfold position_is_final. simpl.
  apply Nat.leb_le. lia.
Qed.

(** * Composition Lemma *)

(** Running on concatenated dictionaries *)
Lemma run_concat : forall alg query n dict1 dict2 s s',
  automaton_run alg query n dict1 s = Some s' ->
  automaton_run alg query n (dict1 ++ dict2) s =
  automaton_run alg query n dict2 s'.
Proof.
  intros alg query n dict1.
  induction dict1 as [| c rest IH]; intros dict2 s s' Hrun.
  - simpl in *. inversion Hrun. subst. reflexivity.
  - simpl in *.
    destruct (transition_state alg s c query n) as [s''|] eqn:Htrans.
    + apply IH. exact Hrun.
    + discriminate.
Qed.

(** * Initial State Properties *)

Lemma initial_state_not_empty : forall alg qlen,
  positions (initial_state alg qlen) <> [].
Proof.
  intros alg qlen.
  unfold initial_state. simpl.
  discriminate.
Qed.

Lemma initial_position_in_initial_state : forall alg qlen,
  In initial_position (positions (initial_state alg qlen)).
Proof.
  intros alg qlen.
  unfold initial_state. simpl.
  left. reflexivity.
Qed.

(** * Examples *)

Example accept_empty_query_empty_dict :
  (* Empty query, empty dict -> distance 0 *)
  forall alg,
  automaton_accepts alg [] 2 [] = true.
Proof.
  intros alg.
  unfold automaton_accepts, automaton_run_from_initial.
  simpl.
  unfold state_is_final, position_is_final. simpl.
  reflexivity.
Qed.

(** Example: Same single-char word should be accepted.
    This would require expanding transition_state which involves
    complex case analysis. Instead, we rely on the soundness/completeness
    theorems which guarantee this property.

    In a full development, this could be proven by:
    1. Computing the actual transition
    2. Showing the final state contains a position (1, 0)
    3. Showing this position is final for query of length 1
*)


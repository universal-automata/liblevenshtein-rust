(** * Levenshtein Distance Core Algorithm

    This module defines the Levenshtein distance function using well-founded
    recursion and provides basic unfolding lemmas.

    Part of: Liblevenshtein.Core

    Decomposed from: Distance.v (lines 62-151)
*)

From Coq Require Import String List Arith Ascii Bool Nat Lia Wf_nat.
From Coq Require Import Program.Wf.
From Coq Require Import Recdef.
Import ListNotations.

From Liblevenshtein.Core Require Import Core.Definitions.

(** * Recursive Definition (Wagner-Fischer Recurrence) *)

(** The Levenshtein distance is defined recursively as the minimum number
    of single-character edits (insertions, deletions, substitutions) needed
    to transform one string into another.

    We use well-founded recursion with measure (length s1 + length s2).
    Each recursive call strictly decreases this measure, guaranteeing termination.
    The Function command generates both the function and proof obligations,
    plus an equation lemma for unfolding. *)

(** Measure function for termination: sum of both string lengths *)
Definition lev_measure (p : list Char * list Char) : nat :=
  length (fst p) + length (snd p).

(** The Levenshtein distance function on pairs, defined using Function
    which provides automatic equation lemmas. Termination is guaranteed
    because each recursive call decreases the total length. *)
Function lev_distance_pair (p : list Char * list Char) {measure lev_measure p} : nat :=
  match p with
  | ([], s2) => length s2
  | (s1, []) => length s1
  | (c1 :: s1', c2 :: s2') =>
      min3 (lev_distance_pair (s1', c2 :: s2') + 1)    (* Delete c1 *)
           (lev_distance_pair (c1 :: s1', s2') + 1)    (* Insert c2 *)
           (lev_distance_pair (s1', s2') + subst_cost c1 c2)  (* Substitute/keep *)
  end.
Proof.
  - (* Termination for diagonal call *)
    intros. unfold lev_measure. simpl. lia.
  - (* Termination for insertion call *)
    intros. unfold lev_measure. simpl. lia.
  - (* Termination for deletion call *)
    intros. unfold lev_measure. simpl. lia.
Defined.

(** Wrapper function with standard signature *)
Definition lev_distance (s1 s2 : list Char) : nat := lev_distance_pair (s1, s2).

(** * Unfolding Lemmas *)

(** Unfolding lemma for lev_distance.
    This follows directly from the equation lemma generated by Function. *)
Lemma lev_distance_unfold : forall s1 s2,
  lev_distance s1 s2 =
    match s1, s2 with
    | [], _ => length s2
    | _, [] => length s1
    | c1 :: s1', c2 :: s2' =>
        min3 (lev_distance s1' s2 + 1)
             (lev_distance s1 s2' + 1)
             (lev_distance s1' s2' + subst_cost c1 c2)
    end.
Proof.
  intros s1 s2.
  unfold lev_distance.
  rewrite lev_distance_pair_equation.
  destruct s1 as [|c1 s1']; [reflexivity|].
  destruct s2 as [|c2 s2']; [reflexivity|].
  reflexivity.
Qed.

(** Base cases for empty strings *)
Lemma lev_distance_empty_left :
  forall s, lev_distance [] s = length s.
Proof.
  intro s.
  rewrite lev_distance_unfold.
  reflexivity.
Qed.

Lemma lev_distance_empty_right :
  forall s, lev_distance s [] = length s.
Proof.
  intro s.
  rewrite lev_distance_unfold.
  destruct s; reflexivity.
Qed.

(** Recursive case *)
Lemma lev_distance_cons :
  forall c1 c2 s1 s2,
    lev_distance (c1 :: s1) (c2 :: s2) =
    min3
      (lev_distance s1 (c2 :: s2) + 1)          (* Delete c1 *)
      (lev_distance (c1 :: s1) s2 + 1)          (* Insert c2 *)
      (lev_distance s1 s2 + subst_cost c1 c2).  (* Substitute/keep *)
Proof.
  intros c1 c2 s1 s2.
  rewrite lev_distance_unfold.
  reflexivity.
Qed.

(** * Position Skipping Optimization - Formal Verification

    This module analyzes the position skipping optimization for sequential rule application.

    **Optimization**: After applying a rule at position `last_pos`, start the next
    iteration's search from `last_pos` instead of position 0.

    **Goal**: Prove whether this optimization preserves semantics or find counterexample.
*)

Require Import String List Arith Ascii Bool Nat Lia.
Require Import PhoneticRewrites.rewrite_rules.
Import ListNotations.

(** * Helper Functions for Optimized Algorithm *)

(** Check if a rule can apply at a position without allocating result *)
Definition can_apply_at (r : RewriteRule) (s : PhoneticString) (pos : nat) : bool :=
  if context_matches (context r) s pos then
    pattern_matches_at (pattern r) s pos
  else
    false.

(** Find first match starting from a given position *)
Fixpoint find_first_match_from (r : RewriteRule) (s : PhoneticString)
                                (start_pos : nat) (remaining : nat) : option nat :=
  match remaining with
  | O => None
  | S remaining' =>
      if can_apply_at r s start_pos then
        Some start_pos
      else
        find_first_match_from r s (S start_pos) remaining'
  end.

(** * Optimized Algorithm *)

(** Sequential rule application with position skipping *)
Fixpoint apply_rules_seq_opt (rules : list RewriteRule) (s : PhoneticString)
                               (fuel : nat) (last_pos : nat)
  : option PhoneticString :=
  match fuel with
  | O => Some s
  | S fuel' =>
      match rules with
      | [] => Some s
      | r :: rest =>
          (** Start search from last_pos instead of 0 *)
          let search_len := (length s - last_pos + 1)%nat in
          match find_first_match_from r s last_pos search_len with
          | Some pos =>
              match apply_rule_at r s pos with
              | Some s' =>
                  (** Rule applied - restart with new last_pos *)
                  apply_rules_seq_opt rules s' fuel' pos
              | None =>
                  (** Shouldn't happen if can_apply_at worked correctly *)
                  apply_rules_seq_opt rest s fuel' last_pos
              end
          | None =>
              (** No match from last_pos onward - try next rule *)
              apply_rules_seq_opt rest s fuel' last_pos
          end
      end
  end.

(** * Key Lemmas *)

(** Lemma: find_first_match_from only searches from start_pos onward *)
Lemma find_first_match_from_lower_bound :
  forall r s start_pos n pos,
    find_first_match_from r s start_pos n = Some pos ->
    (start_pos <= pos)%nat.
Proof.
  intros r s start_pos n.
  generalize dependent start_pos.
  induction n as [| n' IH]; intros start_pos pos H.
  - (* Base case: n = 0 *)
    simpl in H. discriminate H.
  - (* Inductive case *)
    simpl in H.
    destruct (can_apply_at r s start_pos) eqn:E.
    + (* Match found at start_pos *)
      injection H as H_eq.
      subst. lia.
    + (* No match, continue searching *)
      apply IH in H.
      lia.
Qed.

(** Lemma: find_first_match_from with insufficient range returns None *)
Lemma find_first_match_from_empty :
  forall r s start_pos,
    (start_pos > length s)%nat ->
    find_first_match_from r s start_pos 0 = None.
Proof.
  intros. simpl. reflexivity.
Qed.

(** * Termination *)

(** Both algorithms terminate with sufficient fuel *)
Theorem apply_rules_seq_opt_terminates :
  forall rules s fuel last_pos,
    exists result,
      apply_rules_seq_opt rules s fuel last_pos = Some result.
Proof.
  intros rules s fuel last_pos.
  generalize dependent last_pos.
  generalize dependent s.
  generalize dependent rules.
  induction fuel as [| fuel' IH]; intros rules s last_pos.
  - (* Base case: fuel = 0 *)
    exists s.
    simpl. reflexivity.
  - (* Inductive case: fuel = S fuel' *)
    destruct rules as [| r rest].
    + (* No rules *)
      exists s.
      simpl. reflexivity.
    + (* At least one rule *)
      simpl.
      destruct (find_first_match_from r s last_pos (length s - last_pos + 1)) eqn:E_find.
      * (* Match found at position n *)
        destruct (apply_rule_at r s n) eqn:E_apply.
        ** (* Rule applied successfully *)
          (* Recursive call with transformed string *)
          apply (IH (r :: rest) p n).
        ** (* Rule application failed *)
          apply (IH rest s last_pos).
      * (* No match found *)
        apply (IH rest s last_pos).
Qed.

(** * Correctness Analysis *)

(** The key question: when does position skipping preserve semantics? *)

(** If a rule cannot apply at any position < start_pos in the current string,
    then starting the search from start_pos is safe *)
Definition no_early_matches (r : RewriteRule) (s : PhoneticString) (start_pos : nat) : Prop :=
  forall pos, (pos < start_pos)%nat -> can_apply_at r s pos = false.

(** * Auxiliary Lemmas for Arithmetic and Bounds *)

(** Helper lemmas for reasoning about truncating natural number subtraction *)

Lemma sub_add_inverse : forall a b,
  (b <= a)%nat -> (a - b + b = a)%nat.
Proof.
  intros a b H.
  lia.
Qed.

Lemma sub_S_decompose : forall a b,
  (S b <= a)%nat -> (a - S b = a - b - 1)%nat.
Proof.
  intros a b H.
  lia.
Qed.

Lemma sub_lt_mono : forall a b c,
  (a - S b <= c)%nat -> (S b <= a)%nat -> (a - b <= S c)%nat.
Proof.
  intros a b c H H_bound.
  lia.
Qed.

Lemma pos_in_search_range : forall start_pos n pos,
  (pos < start_pos + n)%nat -> (start_pos <= pos)%nat -> (pos - start_pos < n)%nat.
Proof.
  intros start_pos n pos H H_ge.
  lia.
Qed.

Lemma search_range_bound : forall (s : PhoneticString) start_pos pos,
  (pos < start_pos + (length s - start_pos + 1))%nat ->
  (start_pos <= length s)%nat ->
  (pos <= length s)%nat.
Proof.
  intros s start_pos pos H H_bound.
  lia.
Qed.

Lemma search_range_strict_bound : forall (s : PhoneticString) start_pos pos,
  (pos < start_pos + (length s - start_pos + 1))%nat ->
  (start_pos <= length s)%nat ->
  (pos < length s + 1)%nat.
Proof.
  intros s start_pos pos H H_bound.
  assert (H_rewrite: (start_pos + (length s - start_pos + 1) = length s + 1)%nat).
  { lia. }
  rewrite H_rewrite in H.
  exact H.
Qed.

(** * Pattern Non-Emptiness Lemmas *)

(** Well-formed rules have non-empty patterns *)
Lemma pattern_non_empty : forall r,
  wf_rule r -> (length (pattern r) > 0)%nat.
Proof.
  intros r H.
  unfold wf_rule in H.
  destruct H as [H_len H_weight].
  exact H_len.
Qed.

(** Pattern matching requires sufficient space *)
Lemma pattern_matches_at_requires_space : forall pat s pos,
  (length pat > 0)%nat ->
  (pos >= length s)%nat ->
  pattern_matches_at pat s pos = false.
Proof.
  intros pat s pos H_len H_pos.
  destruct pat as [| p ps] eqn:E_pat.
  - (* pat = [], contradicts H_len *)
    simpl in H_len. lia.
  - (* pat = p :: ps, so pattern is non-empty *)
    simpl.
    (* nth_error s pos when pos >= length s returns None *)
    assert (H_nth: nth_error s pos = None).
    { apply nth_error_None. lia. }
    rewrite H_nth.
    reflexivity.
Qed.

(** can_apply_at returns false at or beyond string length for non-empty patterns *)
Lemma can_apply_at_beyond_length : forall r s pos,
  wf_rule r ->
  (pos >= length s)%nat ->
  can_apply_at r s pos = false.
Proof.
  intros r s pos H_wf H_pos.
  unfold can_apply_at.
  destruct (context_matches (context r) s pos) eqn:E_ctx.
  - (* Context matches - check pattern *)
    assert (H_pat_len: (length (pattern r) > 0)%nat).
    { apply pattern_non_empty. exact H_wf. }
    rewrite (pattern_matches_at_requires_space (pattern r) s pos H_pat_len H_pos).
    reflexivity.
  - (* Context doesn't match *)
    reflexivity.
Qed.

(** * Helper Lemmas for Phase 3 *)

(** ** Arithmetic Helpers *)

(** Fuel bound shift: If lower bound holds for fuel, it holds for S fuel *)
Lemma fuel_bound_shift : forall (s : PhoneticString) fuel pos,
  (length s - fuel <= pos)%nat ->
  (length s - S fuel <= pos)%nat.
Proof.
  intros s fuel pos H.
  lia.
Qed.

(** Range arithmetic simplification *)
Lemma range_arithmetic : forall n,
  (n - 0 + 1 = S n)%nat.
Proof.
  intros n.
  lia.
Qed.

(** Natural number subtraction with successor *)
Lemma nat_sub_succ : forall n m,
  (n >= S m)%nat ->
  (n - S m = n - m - 1)%nat.
Proof.
  intros n m H.
  lia.
Qed.

(** ** List Helpers *)

(** Element at head of list *)
Lemma In_head : forall {A : Type} (x : A) (xs : list A),
  In x (x :: xs).
Proof.
  intros A x xs.
  simpl.
  left.
  reflexivity.
Qed.

(** If element in tail, it's in the whole list *)
Lemma In_tail : forall {A : Type} (x y : A) (xs : list A),
  In x xs ->
  In x (y :: xs).
Proof.
  intros A x y xs H.
  simpl.
  right.
  exact H.
Qed.

(** ** Well-formedness Helpers *)

(** Well-formedness preserved for rules in list *)
Lemma wf_rule_In : forall r rules,
  (forall r', In r' rules -> wf_rule r') ->
  In r rules ->
  wf_rule r.
Proof.
  intros r rules H_all H_in.
  apply H_all.
  exact H_in.
Qed.

(** ** Search Helpers *)

(** Generalized can_apply_beyond_length for rules in a list *)
Lemma can_apply_beyond_length_general : forall rules r s pos,
  (forall r', In r' rules -> wf_rule r') ->
  In r rules ->
  (pos >= length s)%nat ->
  can_apply_at r s pos = false.
Proof.
  intros rules r s pos H_wf_all H_in H_pos.
  apply can_apply_at_beyond_length.
  - apply wf_rule_In with (rules := rules); assumption.
  - exact H_pos.
Qed.

(** If apply_rule_at succeeds on a well-formed rule, position must be valid *)
Lemma apply_rule_at_pos_valid : forall r s pos s',
  wf_rule r ->
  apply_rule_at r s pos = Some s' ->
  (pos < length s)%nat.
Proof.
  intros r s pos s' H_wf H_apply.
  (* Proof by contradiction: assume pos >= length s *)
  destruct (lt_dec pos (length s)) as [H_lt | H_ge].
  - (* pos < length s - this is what we want to prove *)
    exact H_lt.
  - (* pos >= length s - show this leads to contradiction *)
    (* If pos >= length s, then apply_rule_at should return None for well-formed rules *)
    unfold apply_rule_at in H_apply.
    destruct (context_matches (context r) s pos) eqn:E_ctx; try discriminate.
    destruct (pattern_matches_at (pattern r) s pos) eqn:E_pat; try discriminate.
    (* But we know pattern_matches_at returns false when pos >= length s for non-empty patterns *)
    assert (H_pat_false: pattern_matches_at (pattern r) s pos = false).
    { apply pattern_matches_at_requires_space.
      - apply pattern_non_empty. exact H_wf.
      - lia. }
    rewrite H_pat_false in E_pat.
    discriminate.
Qed.

(** * Auxiliary Lemmas for find_first_match *)

(** Lemma: find_first_match returns Some only if can_apply_at is true at that position *)
Lemma find_first_match_some_implies_can_apply :
  forall r s fuel pos,
    find_first_match r s fuel = Some pos ->
    can_apply_at r s pos = true.
Proof.
  intros r s fuel.
  generalize dependent s.
  induction fuel as [| fuel' IH]; intros s pos H.
  - (* Base case: fuel = 0 *)
    simpl in H. discriminate H.
  - (* Inductive case *)
    simpl in H.
    unfold is_Some in H.
    destruct (apply_rule_at r s (length s - S fuel')%nat) eqn:E.
    + (* Match found *)
      injection H as H_eq.
      subst pos.
      unfold apply_rule_at in E.
      destruct (context_matches (context r) s (length s - S fuel')%nat) eqn:E_ctx; try discriminate.
      destruct (pattern_matches_at (pattern r) s (length s - S fuel')%nat) eqn:E_pat; try discriminate.
      unfold can_apply_at.
      rewrite E_ctx, E_pat.
      reflexivity.
    + (* No match, continue *)
      apply IH in H.
      exact H.
Qed.

(** Lemma: find_first_match searches from position (length s - fuel) onward *)
Lemma find_first_match_search_range :
  forall r s fuel pos,
    wf_rule r ->
    find_first_match r s fuel = Some pos ->
    (length s - fuel <= pos)%nat /\ (pos < length s)%nat.
Proof.
  intros r s fuel pos H_wf H_match.
  revert s pos H_match.
  induction fuel as [| fuel' IH]; intros s pos H.
  - (* Base case *)
    simpl in H. discriminate H.
  - (* Inductive case *)
    simpl in H.
    destruct (is_Some (apply_rule_at r s (length s - S fuel')%nat)) eqn:E.
    + (* Match found at (length s - S fuel') *)
      injection H as H_eq.
      split.
      * (* Show length s - S fuel' >= length s - fuel' *)
        rewrite <- H_eq. lia.
      * (* Show pos < length s *)
        rewrite <- H_eq.
        (* Position must be < length s *)
        (* When fuel = S fuel', we check position (length s - S fuel') *)
        (* Two cases: either S fuel' <= length s, or S fuel' > length s *)
        destruct (le_lt_dec (S fuel') (length s)) as [H_fuel_bound | H_fuel_large].
        ** (* S fuel' <= length s, so position = length s - S fuel' < length s *)
           lia.
        ** (* S fuel' > length s, so length s - S fuel' = 0 due to truncating subtraction *)
           assert (H_pos_zero: (length s - S fuel' = 0)%nat) by lia.
           rewrite H_pos_zero.
           (* Need to show 0 < length s *)
           (* If apply_rule_at succeeded at position 0, the string must be non-empty *)
           destruct s as [| phone rest] eqn:E_s.
           *** (* s = [], empty string *)
               (* Empty string with apply_rule_at succeeding contradicts well-formedness *)
               (* For well-formed rules, apply_rule_at on empty string at any position returns None *)
               unfold is_Some in E.
               simpl in E.
               (* apply_rule_at r [] 0 with non-empty pattern must be None *)
               assert (H_apply_false: apply_rule_at r [] 0 = None).
               { unfold apply_rule_at.
                 destruct (context_matches (context r) [] 0) eqn:E_ctx.
                 - (* Context matches, but pattern matching on empty string with non-empty pattern fails *)
                   assert (H_pat: pattern_matches_at (pattern r) [] 0 = false).
                   { apply pattern_matches_at_requires_space.
                     - apply pattern_non_empty. exact H_wf.
                     - simpl. lia. }
                   rewrite H_pat. reflexivity.
                 - reflexivity. }
               rewrite H_apply_false in E.
               simpl in E. discriminate E.
           *** (* s = phone :: rest, non-empty *)
               simpl. lia.
    + (* No match, continue *)
      apply (IH s pos) in H.
      destruct H as [H_lower H_upper].
      split; lia.
Qed.

(** Lemma: If find_first_match finds a position, no earlier position matches *)
Lemma find_first_match_is_first :
  forall r s fuel pos,
    find_first_match r s fuel = Some pos ->
    forall p, (p < pos)%nat -> (length s - fuel <= p)%nat -> can_apply_at r s p = false.
Proof.
  intros r s fuel.
  generalize dependent s.
  induction fuel as [| fuel' IH]; intros s pos H p H_less H_ge.
  - (* Base case *)
    simpl in H. discriminate H.
  - (* Inductive case *)
    simpl in H.
    destruct (is_Some (apply_rule_at r s (length s - S fuel')%nat)) eqn:E.
    + (* Match found at (length s - S fuel') *)
      injection H as H_eq.
      subst pos.
      (* p < length s - S fuel', but p >= length s - S fuel', contradiction *)
      assert (H_eq_p: (p = length s - S fuel' \/ p < length s - S fuel')%nat).
      { lia. }
      destruct H_eq_p as [H_eq | H_lt].
      * (* p = length s - S fuel' *)
        subst p.
        lia. (* Contradiction: p < pos but p = pos *)
      * (* p < length s - S fuel' *)
        (* But p >= length s - S fuel', contradiction *)
        lia.
    + (* No match at (length s - S fuel'), continue searching *)
      (* Need to show that can_apply_at at (length s - S fuel') is false *)
      assert (H_range: (length s - S fuel' <= p)%nat /\ (p < pos)%nat).
      { lia. }
      destruct H_range as [H_ge' H_lt'].
      assert (H_eq_or: (p = length s - S fuel' \/ p > length s - S fuel')%nat).
      { lia. }
      destruct H_eq_or as [H_eq | H_gt].
      * (* p = length s - S fuel' *)
        subst p.
        (* apply_rule_at returned None, so can_apply_at must be false *)
        unfold is_Some in E.
        destruct (apply_rule_at r s (length s - S fuel')%nat) eqn:E_apply; try discriminate.
        unfold apply_rule_at in E_apply.
        unfold can_apply_at.
        destruct (context_matches (context r) s (length s - S fuel')%nat) eqn:E_ctx.
        ** (* context matches *)
           destruct (pattern_matches_at (pattern r) s (length s - S fuel')%nat) eqn:E_pat.
           *** (* pattern also matches - but apply_rule_at returned None, contradiction *)
               discriminate E_apply.
           *** (* pattern doesn't match - can_apply_at returns false *)
               reflexivity.
        ** (* context doesn't match - can_apply_at returns false *)
           reflexivity.
      * (* p > length s - S fuel' *)
        apply (IH s pos H p H_lt').
        lia.
Qed.

(** Lemma: If can_apply_at is true at pos and false before, find_first_match finds pos *)
Lemma find_first_match_finds_first_true :
  forall r s fuel pos,
    (pos < length s)%nat ->
    (length s - fuel <= pos)%nat ->
    can_apply_at r s pos = true ->
    (forall p, (length s - fuel <= p)%nat -> (p < pos)%nat -> can_apply_at r s p = false) ->
    find_first_match r s fuel = Some pos.
Proof.
  intros r s fuel pos H_pos_valid H_fuel_bound H_can_apply H_first.

  (* Induction on fuel *)
  induction fuel as [| fuel' IH].
  - (* Base case: fuel = 0 *)
    (* length s - 0 <= pos, so length s <= pos *)
    simpl in H_fuel_bound.
    (* But pos < length s, contradiction *)
    lia.

  - (* Inductive case: fuel = S fuel' *)
    simpl.
    (* Current position: length s - S fuel' *)
    destruct (Nat.eq_dec pos (length s - S fuel')) as [H_pos_eq | H_pos_ne].

    + (* Case 1: pos = length s - S fuel', we should find it immediately *)
      subst pos.
      (* is_Some (apply_rule_at ...) = true because can_apply_at is true *)
      assert (H_is_some_true: is_Some (apply_rule_at r s (length s - S fuel')%nat) = true).
      { unfold is_Some.
        unfold apply_rule_at.
        unfold can_apply_at in H_can_apply.
        destruct (context_matches (context r) s (length s - S fuel')%nat) eqn:E_ctx;
        destruct (pattern_matches_at (pattern r) s (length s - S fuel')%nat) eqn:E_pat;
        try discriminate H_can_apply.
        reflexivity. }
      rewrite H_is_some_true.
      reflexivity.

    + (* Case 2: pos ≠ length s - S fuel' *)
      (* Since length s - S fuel' <= pos (from H_fuel_bound) and pos ≠ length s - S fuel',
         we have length s - S fuel' < pos *)
      assert (H_pos_gt: (length s - S fuel' < pos)%nat).
      { lia. }

      (* The current position (length s - S fuel') is in the range and < pos,
         so by H_first, can_apply_at must be false there *)
      assert (H_current_false: can_apply_at r s (length s - S fuel')%nat = false).
      { apply H_first.
        - (* Show length s - S fuel' >= length s - S fuel' *)
          lia.
        - (* Show length s - S fuel' < pos *)
          exact H_pos_gt. }

      (* is_Some (apply_rule_at ...) = false when can_apply_at is false *)
      assert (H_is_some_false: is_Some (apply_rule_at r s (length s - S fuel')%nat) = false).
      { unfold is_Some, apply_rule_at.
        unfold can_apply_at in H_current_false.
        destruct (context_matches (context r) s (length s - S fuel')%nat) eqn:E_ctx.
        - (* context matches *)
          simpl in H_current_false.
          destruct (pattern_matches_at (pattern r) s (length s - S fuel')%nat) eqn:E_pat.
          + (* pattern matches - contradiction *)
            discriminate H_current_false.
          + (* pattern doesn't match *)
            reflexivity.
        - (* context doesn't match *)
          reflexivity. }

      rewrite H_is_some_false.

      (* Use IH on fuel' *)
      apply IH.
      * (* Show length s - fuel' <= pos *)
        (* We have length s - S fuel' < pos from H_pos_gt *)
        (* length s - fuel' = length s - S fuel' + 1 when non-truncating *)
        (* So length s - S fuel' < pos implies length s - fuel' <= pos *)
        destruct (le_lt_dec (S fuel') (length s)) as [H_fuel_ok | H_fuel_large].
        ** (* S fuel' <= length s, non-truncating case *)
           (* length s - fuel' = (length s - S fuel') + 1 *)
           (* Since length s - S fuel' < pos, we have (length s - S fuel') + 1 <= pos *)
           lia.
        ** (* S fuel' > length s, both truncate to 0 *)
           assert (H_zero: (length s - fuel' = 0)%nat) by lia.
           rewrite H_zero.
           lia.
      * (* Show all positions in [length s - fuel', pos) have can_apply_at false *)
        intros p H_p_ge H_p_lt.
        apply H_first.
        ** (* Show length s - S fuel' <= p *)
           (* We have length s - fuel' <= p *)
           (* Since S fuel' > fuel', we have length s - S fuel' < length s - fuel' *)
           (* Therefore length s - S fuel' <= p *)
           transitivity (length s - fuel')%nat.
           *** (* length s - S fuel' <= length s - fuel' *)
               destruct (le_lt_dec (S fuel') (length s)) as [H_fuel_ok | H_fuel_large].
               **** lia.
               **** (* S fuel' > length s, both sides truncate to 0 *)
                    assert (H1: (length s - S fuel' = 0)%nat) by lia.
                    assert (H2: (length s - fuel' = 0)%nat) by lia.
                    rewrite H1, H2. lia.
           *** exact H_p_ge.
        ** exact H_p_lt.
Qed.

(** Lemma: find_first_match_from returns positions within bounds *)
Lemma find_first_match_from_upper_bound :
  forall r s start_pos n pos,
    find_first_match_from r s start_pos n = Some pos ->
    (pos < start_pos + n)%nat.
Proof.
  intros r s start_pos n.
  generalize dependent start_pos.
  induction n as [| n' IH]; intros start_pos pos H.
  - simpl in H. discriminate.
  - simpl in H.
    destruct (can_apply_at r s start_pos) eqn:E.
    + injection H as H_eq. subst. lia.
    + apply IH in H. lia.
Qed.

(** Lemma: find_first_match_from is "first" - no earlier position matches *)
Lemma find_first_match_from_is_first :
  forall r s start_pos n pos,
    find_first_match_from r s start_pos n = Some pos ->
    forall p, (start_pos <= p)%nat -> (p < pos)%nat -> can_apply_at r s p = false.
Proof.
  intros r s start_pos n.
  generalize dependent start_pos.
  induction n as [| n' IH]; intros start_pos pos H p H_ge H_lt.
  - simpl in H. discriminate.
  - simpl in H.
    destruct (can_apply_at r s start_pos) eqn:E.
    + (* Match found at start_pos *)
      injection H as H_eq. subst.
      (* p < pos = start_pos, but p >= start_pos, contradiction *)
      lia.
    + (* No match at start_pos, continue *)
      assert (H_eq_or: (p = start_pos \/ p > start_pos)%nat).
      { lia. }
      destruct H_eq_or as [H_eq | H_gt].
      * subst. exact E.
      * apply (IH (S start_pos) pos H p); lia.
Qed.

(** Helper: find_first_match_from returns positions where can_apply_at is true *)
Lemma find_first_match_from_implies_can_apply :
  forall r s start_pos n pos,
    find_first_match_from r s start_pos n = Some pos ->
    can_apply_at r s pos = true.
Proof.
  intros r s start_pos n.
  generalize dependent start_pos.
  induction n as [| n' IH]; intros start_pos pos H.
  - (* Base case: n = 0 *)
    simpl in H. discriminate.
  - (* Inductive case *)
    simpl in H.
    destruct (can_apply_at r s start_pos) eqn:E.
    + (* Found match at start_pos *)
      injection H as H_eq. subst. exact E.
    + (* Continue search *)
      apply (IH (S start_pos) pos H).
Qed.

(** Generalized equivalence lemma with arbitrary fuel and start position *)
Lemma find_first_match_equiv_general :
  forall r s fuel start_pos,
    wf_rule r ->
    start_pos = (length s - fuel)%nat ->
    (fuel <= length s)%nat ->
    find_first_match r s fuel = find_first_match_from r s start_pos (fuel + 1)%nat.
Proof.
  intros r s fuel start_pos H_wf H_start H_fuel_bound.
  subst start_pos.

  (* Induction on fuel *)
  induction fuel as [| fuel' IH].

  - (* Base case: fuel = 0 *)
    simpl.
    (* LHS: None *)
    (* RHS: find_first_match_from r s (length s) 1 *)
    assert (H_zero: (length s - 0 = length s)%nat) by lia.
    rewrite H_zero.
    simpl.
    (* Position length s is out of bounds, so can_apply_at returns false *)
    assert (H_out_of_bounds: can_apply_at r s (length s) = false).
    { apply can_apply_at_beyond_length; try assumption. lia. }
    rewrite H_out_of_bounds.
    reflexivity.

  - (* Inductive case: fuel = S fuel' *)
    simpl.
    (* Both check position (length s - S fuel') *)
    (* Note: S fuel' + 1 simplifies to S (S fuel') *)

    (* Case split on whether rule applies at current position *)
    destruct (can_apply_at r s (length s - S fuel')%nat) eqn:E_apply.

    + (* Rule applies at current position *)
      (* LHS: is_Some (apply_rule_at ...) should be true *)
      unfold is_Some, apply_rule_at, can_apply_at in *.
      destruct (context_matches (context r) s (length s - S fuel')%nat) eqn:E_ctx;
      destruct (pattern_matches_at (pattern r) s (length s - S fuel')%nat) eqn:E_pat;
      try discriminate E_apply.
      reflexivity.

    + (* Rule doesn't apply at current position *)
      (* LHS: is_Some (apply_rule_at ...) should be false *)
      (* RHS: find_first_match_from recurses *)
      unfold is_Some, apply_rule_at in *.
      unfold can_apply_at in E_apply.

      (* Both functions recurse to next position *)
      (* Need to relate: find_first_match r s fuel'
                    and: find_first_match_from r s (S (length s - S fuel')) (S fuel') *)

      (* Show S (length s - S fuel') = length s - fuel' *)
      assert (H_pos_shift: (S (length s - S fuel') = length s - fuel')%nat).
      { destruct (le_lt_dec (S fuel') (length s)) as [H_ok | H_large].
        - lia.
        - (* S fuel' > length s contradicts H_fuel_bound *)
          lia. }

      (* Rewrite based on can_apply_at being false *)
      destruct (context_matches (context r) s (length s - S fuel')%nat) eqn:E_ctx.
      * (* Context matches but pattern doesn't *)
        destruct (pattern_matches_at (pattern r) s (length s - S fuel')%nat) eqn:E_pat.
        ** (* Both true - contradiction with E_apply *)
           simpl in E_apply. discriminate E_apply.
        ** (* Context true, pattern false *)
           rewrite H_pos_shift.
           rewrite IH; try lia.
           reflexivity.
      * (* Context doesn't match *)
        rewrite H_pos_shift.
        rewrite IH; try lia.
        reflexivity.
Qed.

(** Lemma: find_first_match and find_first_match_from starting at 0 are equivalent *)
Lemma find_first_match_equiv_from_zero :
  forall r s,
    wf_rule r ->
    find_first_match r s (length s) = find_first_match_from r s 0 (length s - 0 + 1)%nat.
Proof.
  intros r s H_wf.
  (* Simplify: length s - 0 + 1 = S (length s) *)
  assert (H_simpl: (length s - 0 + 1 = S (length s))%nat) by lia.
  rewrite H_simpl.

  (* Use generalized equivalence with fuel = length s *)
  (* Note: length s - length s = 0, and length s + 1 = S (length s) *)
  assert (H_eq: find_first_match r s (length s) =
                find_first_match_from r s (length s - length s)%nat (length s + 1)%nat).
  { apply find_first_match_equiv_general; try assumption.
    - reflexivity.
    - lia. }

  (* Simplify: length s - length s = 0, length s + 1 = S (length s) *)
  assert (H_zero: (length s - length s = 0)%nat) by lia.
  assert (H_succ: (length s + 1 = S (length s))%nat) by lia.
  rewrite H_zero, H_succ in H_eq.
  exact H_eq.
Qed.

(** Lemma: Reverse direction - from find_first_match_from to find_first_match *)
Lemma find_first_match_equiv_from_zero_reverse :
  forall r s pos,
    wf_rule r ->
    find_first_match_from r s 0 (length s - 0 + 1)%nat = Some pos ->
    find_first_match r s (length s) = Some pos.
Proof.
  intros r s pos H_wf H_from.
  assert (H_equiv: find_first_match r s (length s) =
                   find_first_match_from r s 0 (length s - 0 + 1)%nat).
  { apply find_first_match_equiv_from_zero. exact H_wf. }
  rewrite H_equiv.
  exact H_from.
Qed.

(** Lemma: Bidirectional equivalence between find_first_match and find_first_match_from from 0 *)
Lemma find_first_match_from_zero_bidirectional :
  forall r s,
    wf_rule r ->
    find_first_match r s (length s) = find_first_match_from r s 0 (length s - 0 + 1)%nat.
Proof.
  intros r s H_wf.
  apply find_first_match_equiv_from_zero.
  exact H_wf.
Qed.

(** * Position-Independence Infrastructure *)

(** Lemma: apply_rule_at preserves phones before the match position *)
Lemma apply_rule_at_preserves_prefix :
  forall r s pos s',
    wf_rule r ->
    apply_rule_at r s pos = Some s' ->
    (forall i, (i < pos)%nat -> nth_error s i = nth_error s' i).
Proof.
  intros r s pos s' H_wf H_apply i H_lt.

  (* First, establish that pos < length s using existing lemma *)
  assert (H_pos_valid: (pos < length s)%nat).
  { eapply apply_rule_at_pos_valid; eauto. }

  unfold apply_rule_at in H_apply.
  destruct (context_matches (context r) s pos) eqn:E_ctx; try discriminate.
  destruct (pattern_matches_at (pattern r) s pos) eqn:E_pat; try discriminate.
  injection H_apply as H_s'.

  (* Goal: nth_error s i = nth_error s' i *)
  (* Strategy: Prove each direction separately then combine *)

  (* First, show what nth_error (firstn pos s) i equals *)
  assert (H_firstn_eq: nth_error (firstn pos s) i = nth_error s i).
  {
    rewrite nth_error_firstn.
    (* This gives: if i <? pos then nth_error s i else None *)
    assert (H_ltb: (i <? pos)%nat = true) by (apply Nat.ltb_lt; exact H_lt).
    rewrite H_ltb.
    reflexivity.
  }

  (* Second, show what nth_error s' i equals *)
  assert (H_s'_eq: nth_error s' i = nth_error (firstn pos s) i).
  {
    rewrite <- H_s'.
    (* Goal: nth_error ((firstn pos s) ++ ...) i = nth_error (firstn pos s) i *)
    rewrite nth_error_app1.
    - reflexivity.
    - (* Show i < length (firstn pos s) *)
      rewrite firstn_length.
      rewrite Nat.min_l by lia.
      exact H_lt.
  }

  (* Combine the two *)
  rewrite H_s'_eq.
  rewrite H_firstn_eq.
  reflexivity.
Qed.

(** Definition: A context preserves its truth value at earlier positions after a transformation *)
Definition context_preserved_at_earlier_positions (ctx : Context) (s s' : PhoneticString) (transform_pos : nat) : Prop :=
  forall pos, (pos < transform_pos)%nat ->
    context_matches ctx s pos = context_matches ctx s' pos.

(** Lemma: Initial context is always preserved (only depends on pos = 0) *)
Lemma initial_context_preserved :
  forall s s' transform_pos,
    (transform_pos > 0)%nat ->
    context_preserved_at_earlier_positions Initial s s' transform_pos.
Proof.
  intros s s' transform_pos H_pos_gt.
  unfold context_preserved_at_earlier_positions.
  intros pos H_lt.
  (* Initial only matches at position 0 *)
  unfold context_matches.
  destruct (Nat.eq_dec pos 0) as [H_eq | H_ne].
  - (* pos = 0, and transform_pos > 0, so position 0 is unchanged *)
    subst pos.
    reflexivity.
  - (* pos <> 0, so Initial doesn't match in either case *)
    reflexivity.
Qed.

(** Lemma: Anywhere context is always preserved (always matches) *)
Lemma anywhere_context_preserved :
  forall s s' transform_pos,
    context_preserved_at_earlier_positions Anywhere s s' transform_pos.
Proof.
  intros s s' transform_pos.
  unfold context_preserved_at_earlier_positions.
  intros pos H_lt.
  unfold context_matches.
  reflexivity.
Qed.

(** Lemma: BeforeVowel context is preserved at earlier positions *)
Lemma before_vowel_context_preserved :
  forall vowels s s' transform_pos,
    (forall i, (i < transform_pos)%nat -> nth_error s i = nth_error s' i) ->
    context_preserved_at_earlier_positions (BeforeVowel vowels) s s' transform_pos.
Proof.
  intros vowels s s' transform_pos H_prefix.
  unfold context_preserved_at_earlier_positions.
  intros pos H_lt.
  unfold context_matches.
  (* BeforeVowel checks nth_error s pos *)
  (* We need to show: (match nth_error s pos with ...) = (match nth_error s' pos with ...) *)
  rewrite <- (H_prefix pos H_lt).
  reflexivity.
Qed.

(** Lemma: BeforeConsonant context is preserved at earlier positions *)
Lemma before_consonant_context_preserved :
  forall consonants s s' transform_pos,
    (forall i, (i < transform_pos)%nat -> nth_error s i = nth_error s' i) ->
    context_preserved_at_earlier_positions (BeforeConsonant consonants) s s' transform_pos.
Proof.
  intros consonants s s' transform_pos H_prefix.
  unfold context_preserved_at_earlier_positions.
  intros pos H_lt.
  unfold context_matches.
  (* BeforeConsonant checks nth_error s pos *)
  rewrite <- (H_prefix pos H_lt).
  reflexivity.
Qed.

(** Lemma: AfterConsonant context is preserved at earlier positions *)
Lemma after_consonant_context_preserved :
  forall consonants s s' transform_pos,
    (forall i, (i < transform_pos)%nat -> nth_error s i = nth_error s' i) ->
    context_preserved_at_earlier_positions (AfterConsonant consonants) s s' transform_pos.
Proof.
  intros consonants s s' transform_pos H_prefix.
  unfold context_preserved_at_earlier_positions.
  intros pos H_lt.
  unfold context_matches.
  (* AfterConsonant checks nth_error s (pos - 1) when pos > 0 *)
  destruct pos as [| pos'].
  - (* pos = 0: AfterConsonant returns false in both cases *)
    reflexivity.
  - (* pos = S pos': need to show nth_error s pos' = nth_error s' pos' *)
    assert (H_pos'_lt: (pos' < transform_pos)%nat) by lia.
    rewrite <- (H_prefix pos' H_pos'_lt).
    reflexivity.
Qed.

(** Lemma: AfterVowel context is preserved at earlier positions *)
Lemma after_vowel_context_preserved :
  forall vowels s s' transform_pos,
    (forall i, (i < transform_pos)%nat -> nth_error s i = nth_error s' i) ->
    context_preserved_at_earlier_positions (AfterVowel vowels) s s' transform_pos.
Proof.
  intros vowels s s' transform_pos H_prefix.
  unfold context_preserved_at_earlier_positions.
  intros pos H_lt.
  unfold context_matches.
  (* AfterVowel checks nth_error s (pos - 1) when pos > 0 *)
  destruct pos as [| pos'].
  - (* pos = 0: AfterVowel returns false in both cases *)
    reflexivity.
  - (* pos = S pos': need to show nth_error s pos' = nth_error s' pos' *)
    assert (H_pos'_lt: (pos' < transform_pos)%nat) by lia.
    rewrite <- (H_prefix pos' H_pos'_lt).
    reflexivity.
Qed.

(** * Context Position-Dependence *)

(** A context is position-dependent if it can change truth value when string changes *)
Definition position_dependent_context (ctx : Context) : bool :=
  match ctx with
  | Final => true  (* Depends on string length *)
  | Initial => false  (* Position 0 is invariant *)
  | BeforeVowel _ => false  (* Depends only on local structure *)
  | AfterConsonant _ => false
  | BeforeConsonant _ => false
  | AfterVowel _ => false
  | Anywhere => false
  end.

(** Lemma: Pattern matching is preserved at positions before transformation *)
Lemma pattern_matches_preserved_before_transformation :
  forall pat s s' pos transform_pos,
    (forall i, (i < transform_pos)%nat -> nth_error s i = nth_error s' i) ->
    (pos + length pat <= transform_pos)%nat ->
    pattern_matches_at pat s pos = pattern_matches_at pat s' pos.
Proof.
  intros pat.
  induction pat as [| p ps IH]; intros s s' pos transform_pos H_prefix H_bound.
  - (* Base case: empty pattern *)
    simpl. reflexivity.
  - (* Inductive case: p :: ps *)
    simpl.
    simpl in H_bound.
    (* Check if pos < transform_pos *)
    assert (H_pos_lt: (pos < transform_pos)%nat) by lia.
    (* Rewrite nth_error s pos to nth_error s' pos *)
    rewrite <- (H_prefix pos H_pos_lt).
    destruct (nth_error s pos) as [p'|] eqn:E_nth.
    + (* Phone found at position pos *)
      destruct (Phone_eqb p p') eqn:E_eq.
      * (* Phones match, check rest of pattern *)
        (* Need to show pattern_matches_at ps s (S pos) = pattern_matches_at ps s' (S pos) *)
        apply (IH s s' (S pos) transform_pos).
        ** exact H_prefix.
        ** lia.
      * (* Phones don't match *)
        reflexivity.
    + (* No phone at position pos *)
      reflexivity.
Qed.

(** Lemma: After applying a position-independent rule at pos, no new matches appear before pos
    (for patterns that don't extend into the modified region) *)
Lemma no_new_early_matches_after_transformation :
  forall r s pos s' r' p,
    wf_rule r ->
    wf_rule r' ->
    position_dependent_context (context r') = false ->
    apply_rule_at r s pos = Some s' ->
    (p < pos)%nat ->
    (p + length (pattern r') <= pos)%nat ->  (* Pattern doesn't extend beyond transformation point *)
    can_apply_at r' s' p = true ->
    can_apply_at r' s p = true.
Proof.
  intros r s pos s' r' p H_wf H_wf' H_indep H_apply H_p_lt H_pattern_bound H_can_s'.

  (* Step 1: Extract prefix preservation *)
  assert (H_prefix: forall i, (i < pos)%nat -> nth_error s i = nth_error s' i).
  { intros i H_i_lt.
    apply (apply_rule_at_preserves_prefix r s pos s' H_wf H_apply i H_i_lt).
  }

  (* Step 2: Unfold can_apply_at and analyze H_can_s' *)
  unfold can_apply_at in H_can_s'.
  destruct (context_matches (context r') s' p) eqn:E_ctx_s'; try discriminate.
  destruct (pattern_matches_at (pattern r') s' p) eqn:E_pat_s'; try discriminate.
  clear H_can_s'.

  (* Step 3: Case analysis on context type *)
  unfold can_apply_at.
  destruct (context r') eqn:E_ctx.

  - (* Initial *)
    (* Use context preservation to relate s and s' *)
    assert (H_ctx_eq: context_matches Initial s p = context_matches Initial s' p).
    { pose proof (initial_context_preserved s s' pos) as H_pres.
      assert (H_pos_gt: (pos > 0)%nat) by lia.
      specialize (H_pres H_pos_gt p H_p_lt).
      exact H_pres.
    }
    rewrite H_ctx_eq, E_ctx_s'.
    rewrite (pattern_matches_preserved_before_transformation (pattern r') s s' p pos); auto.



  - (* Final - contradiction *)
    simpl in H_indep.
    discriminate H_indep.

  - (* BeforeVowel *)
    assert (H_ctx_eq: context_matches (BeforeVowel l) s p = context_matches (BeforeVowel l) s' p).
    { pose proof (before_vowel_context_preserved l s s' pos H_prefix p H_p_lt) as H_pres.
      exact H_pres.
    }
    rewrite H_ctx_eq, E_ctx_s'.
    rewrite (pattern_matches_preserved_before_transformation (pattern r') s s' p pos); auto.

  - (* AfterConsonant *)
    assert (H_ctx_eq: context_matches (AfterConsonant l) s p = context_matches (AfterConsonant l) s' p).
    { pose proof (after_consonant_context_preserved l s s' pos H_prefix p H_p_lt) as H_pres.
      exact H_pres.
    }
    rewrite H_ctx_eq, E_ctx_s'.
    rewrite (pattern_matches_preserved_before_transformation (pattern r') s s' p pos); auto.

  - (* BeforeConsonant *)
    assert (H_ctx_eq: context_matches (BeforeConsonant l) s p = context_matches (BeforeConsonant l) s' p).
    { pose proof (before_consonant_context_preserved l s s' pos H_prefix p H_p_lt) as H_pres.
      exact H_pres.
    }
    rewrite H_ctx_eq, E_ctx_s'.
    rewrite (pattern_matches_preserved_before_transformation (pattern r') s s' p pos); auto.

  - (* AfterVowel *)
    assert (H_ctx_eq: context_matches (AfterVowel l) s p = context_matches (AfterVowel l) s' p).
    { pose proof (after_vowel_context_preserved l s s' pos H_prefix p H_p_lt) as H_pres.
      exact H_pres.
    }
    rewrite H_ctx_eq, E_ctx_s'.
    rewrite (pattern_matches_preserved_before_transformation (pattern r') s s' p pos); auto.

  - (* Anywhere *)
    assert (H_ctx_eq: context_matches Anywhere s p = context_matches Anywhere s' p).
    { pose proof (anywhere_context_preserved s s' pos) as H_pres.
      unfold context_preserved_at_earlier_positions in H_pres.
      apply (H_pres p H_p_lt).
    }
    rewrite H_ctx_eq, E_ctx_s'.
    rewrite (pattern_matches_preserved_before_transformation (pattern r') s s' p pos); auto.
Qed.


(** Lemma: If no early matches exist, both find the same match (or both find none) *)
Lemma find_first_match_from_equivalent_when_no_early_matches :
  forall r s start_pos,
    wf_rule r ->
    no_early_matches r s start_pos ->
    (forall pos, find_first_match_from r s start_pos (length s - start_pos + 1) = Some pos ->
                 find_first_match r s (length s) = Some pos).
Proof.
  intros r s start_pos H_wf H_no_early pos H_found.
  unfold no_early_matches in H_no_early.

  (* find_first_match_from found pos, so can_apply_at r s pos = true *)
  assert (H_can_apply: can_apply_at r s pos = true).
  {
    eapply find_first_match_from_implies_can_apply. eauto.
  }

  (* pos >= start_pos *)
  assert (H_bound: (start_pos <= pos)%nat).
  { eapply find_first_match_from_lower_bound. eauto. }

  (* pos < length s: from the search bounds and can_apply_at being true *)
  assert (H_pos_in_bounds: (pos < length s)%nat).
  {
    (* find_first_match_from searched up to position start_pos + n - 1 where n = length s - start_pos + 1 *)
    assert (H_upper: (pos < start_pos + (length s - start_pos + 1))%nat).
    { eapply find_first_match_from_upper_bound. eauto. }
    (* Simplify the bound *)
    destruct (le_lt_dec start_pos (length s)) as [H_start_ok | H_start_large].
    - (* start_pos <= length s, so expression simplifies *)
      assert (H_rewrite: (start_pos + (length s - start_pos + 1) = length s + 1)%nat) by lia.
      rewrite H_rewrite in H_upper.
      (* pos < length s + 1 means pos <= length s *)
      (* To show pos < length s, need to exclude pos = length s *)
      destruct (Nat.eq_dec pos (length s)) as [H_eq | H_ne].
      * (* pos = length s - but can_apply_at at or beyond length s is false for wf rules *)
        subst pos.
        (* This contradicts H_can_apply *)
        assert (H_false: can_apply_at r s (length s) = false).
        { apply can_apply_at_beyond_length. exact H_wf. lia. }
        rewrite H_false in H_can_apply.
        discriminate.
      * (* pos <> length s, and pos <= length s, so pos < length s *)
        lia.
    - (* start_pos > length s, then length s - start_pos = 0 *)
      (* So search range is [start_pos, start_pos + 1) *)
      (* But if can_apply_at is true at pos, and pos >= start_pos > length s *)
      (* This contradicts can_apply_at requiring valid position *)
      (* can_apply_at checks context and pattern at position pos *)
      (* For position >= length s, context matching could succeed, but pattern matching *)
      (* requires pos + pattern_length <= length s, which fails if pos >= length s and pattern non-empty *)
      (* H_upper: pos < start_pos + (length s - start_pos + 1) *)
      (* With length s - start_pos = 0, this becomes pos < start_pos + 1 *)
      (* Which means pos <= start_pos *)
      (* Since start_pos > length s and pos >= start_pos, we have pos >= length s *)
      (* But can_apply_at at position >= length s should be false for non-empty patterns *)
      (* This is getting complex - for now, use a simpler bound *)
      (* Actually, from H_upper, pos < start_pos + 1, so pos <= start_pos *)
      (* Combined with H_bound (start_pos <= pos), we get pos = start_pos *)
      assert (H_pos_eq: pos = start_pos) by lia.
      subst pos.
      (* Now start_pos > length s, but can_apply_at r s start_pos = true *)
      (* This contradicts can_apply_at being false beyond string length for wf rules *)
      assert (H_false: can_apply_at r s start_pos = false).
      { apply can_apply_at_beyond_length. exact H_wf. lia. }
      rewrite H_false in H_can_apply.
      discriminate.
  }

  (* Use find_first_match_finds_first_true to show find_first_match finds pos *)
  apply find_first_match_finds_first_true.
  - exact H_pos_in_bounds.
  - lia.
  - exact H_can_apply.
  - (* For all p in [0, pos), can_apply_at r s p = false *)
    intros p H_range H_lt.
    destruct (Nat.lt_ge_cases p start_pos) as [H_before_start | H_after_start].
    + (* p < start_pos: use H_no_early *)
      apply H_no_early. exact H_before_start.
    + (* start_pos <= p < pos *)
      (* Use find_first_match_from_is_first *)
      eapply find_first_match_from_is_first; eauto.
Qed.

(** * Context-Specific Safety *)

(** Helper Lemma: Skipping a single non-matching position *)
Lemma find_first_match_from_skip_one :
  forall r s pos n,
    can_apply_at r s pos = false ->
    find_first_match_from r s pos (S n) =
    find_first_match_from r s (S pos) n.
Proof.
  intros r s pos n H_no_match.
  simpl.
  rewrite H_no_match.
  reflexivity.
Qed.

(** Helper Lemma: General version - skip from any starting position to any target *)
Lemma find_first_match_from_skip_range :
  forall r s start_from end_at remaining,
    (forall p, (start_from <= p < end_at)%nat -> can_apply_at r s p = false) ->
    (end_at + remaining <= S (length s))%nat ->
    (start_from <= end_at)%nat ->
    find_first_match_from r s start_from (end_at - start_from + remaining) =
    find_first_match_from r s end_at remaining.
Proof.
  intros r s start_from end_at.
  (* Induct on the gap: end_at - start_from *)
  remember (end_at - start_from)%nat as gap.
  revert start_from end_at Heqgap.
  induction gap as [| k IH]; intros start_from end_at Heqgap remaining H_no_match H_bound H_order.

  - (* Base: gap = 0, so start_from = end_at *)
    assert (start_from = end_at) by lia.
    subst.
    replace (end_at - end_at + remaining)%nat with remaining by lia.
    reflexivity.

  - (* Inductive: gap = S k *)
    (* start_from < end_at, so position start_from exists and doesn't match *)
    assert (H_start_no_match: can_apply_at r s start_from = false).
    { apply H_no_match. lia. }

    (* From Heqgap, we know end_at - start_from = S k *)
    (* So the goal's count is: S k + remaining *)

    (* Unfold find_first_match_from once to expose the recursion *)
    destruct (end_at - start_from + remaining)%nat eqn:Hcount.
    + (* Count is 0 - impossible since it equals S k + remaining *)
      exfalso. lia.

    + (* Count is S n0 *)
      simpl.
      rewrite H_start_no_match.

      (* After skipping start_from, we recurse from S start_from with count n0 *)
      (* Apply IH to finish *)
      apply (IH (S start_from) end_at).
      * (* Gap: end_at - S start_from = k *) lia.
      * (* Positions in [S start_from, end_at) don't match *)
        intros p H_p_range.
        apply H_no_match. lia.
      * (* Bound *) lia.
      * (* Order *) lia.
Qed.

(** * Multi-Rule Invariant: Infrastructure for Proving Position-Skipping Safety *)

(** ** Invariant Predicate Definitions *)

(** The fundamental invariant: no rules in the list match at any position before max_pos *)
Definition no_rules_match_before (rules : list RewriteRule) (s : PhoneticString) (max_pos : nat) : Prop :=
  forall r, In r rules -> forall p, (p < max_pos)%nat -> can_apply_at r s p = false.

(** Variant with pattern length constraint: only positions where patterns fit *)
Definition no_rules_match_before_with_space (rules : list RewriteRule) (s : PhoneticString) (max_pos : nat) : Prop :=
  forall r, In r rules ->
    forall p, (p < max_pos)%nat ->
      (p + length (pattern r) <= max_pos)%nat ->
      can_apply_at r s p = false.

(** ** Establishment Lemmas: find_first_match establishes the invariant *)

(** Lemma: When find_first_match finds a position for a single rule,
    all earlier positions don't match *)
Lemma find_first_match_establishes_invariant_single :
  forall r s pos,
    wf_rule r ->
    find_first_match r s (length s) = Some pos ->
    no_rules_match_before [r] s pos.
Proof.
  intros r s pos H_wf H_find.
  unfold no_rules_match_before.
  intros r0 H_in p H_p_lt.
  (* r0 must be r since [r] is a singleton list *)
  destruct H_in as [H_eq | H_in_empty].
  - (* r0 = r *)
    subst r0.
    (* Use find_first_match_is_first lemma *)
    eapply find_first_match_is_first; eauto.
    (* Need to show: length s - length s <= p *)
    lia.
  - (* r0 ∈ [] - impossible *)
    inversion H_in_empty.
Qed.

(** Lemma: The invariant holds for the empty rule list (vacuously true) *)
Lemma no_rules_match_before_empty :
  forall s pos,
    no_rules_match_before [] s pos.
Proof.
  intros s pos.
  unfold no_rules_match_before.
  intros r H_in.
  inversion H_in.  (* No rules in empty list *)
Qed.

(** ** Preservation Lemmas: The invariant is preserved by transformation *)

(** Lemma: If a single rule doesn't match before pos in s,
    it won't match after transformation to s' (with pattern bound constraint) *)
Lemma single_rule_no_match_preserved :
  forall r r_applied s pos s' p,
    wf_rule r_applied ->
    wf_rule r ->
    position_dependent_context (context r) = false ->
    apply_rule_at r_applied s pos = Some s' ->
    (p < pos)%nat ->
    (p + length (pattern r) <= pos)%nat ->  (* Pattern fits before transformation point *)
    can_apply_at r s p = false ->
    can_apply_at r s' p = false.
Proof.
  intros r r_applied s pos s' p H_wf_applied H_wf H_indep H_apply H_p_lt H_pattern_bound H_no_match_s.
  (* Proof by contrapositive of no_new_early_matches_after_transformation *)
  destruct (can_apply_at r s' p) eqn:E_match_s'; try reflexivity.
  (* If can_apply_at r s' p = true, then by no_new_early_matches, can_apply_at r s p = true *)
  assert (H_match_s: can_apply_at r s p = true).
  { apply (no_new_early_matches_after_transformation r_applied s pos s' r p H_wf_applied H_wf H_indep H_apply H_p_lt H_pattern_bound E_match_s'). }
  (* But this contradicts H_no_match_s *)
  rewrite H_match_s in H_no_match_s.
  discriminate H_no_match_s.
Qed.

(** Lemma: If no rules in a list match before pos in s,
    and patterns all fit, then no rules match after transformation *)
Lemma all_rules_no_match_preserved :
  forall rules r_applied s pos s' p,
    wf_rule r_applied ->
    (forall r0, In r0 rules -> wf_rule r0) ->
    (forall r0, In r0 rules -> position_dependent_context (context r0) = false) ->
    (forall r0, In r0 rules -> (p + length (pattern r0) <= pos)%nat) ->  (* All patterns fit *)
    apply_rule_at r_applied s pos = Some s' ->
    (p < pos)%nat ->
    no_rules_match_before rules s pos ->
    no_rules_match_before rules s' p.
Proof.
  intros rules r_applied s pos s' p H_wf_applied H_wf_all H_indep_all H_pattern_bounds H_apply H_p_lt H_inv_before.
  unfold no_rules_match_before in *.
  intros r0 H_in_r0 p0 H_p0_lt.

  (* Get the hypothesis that r0 doesn't match in s *)
  assert (H_r0_no_match_s: can_apply_at r0 s p0 = false).
  { apply H_inv_before.
    - exact H_in_r0.
    - (* p0 < p < pos, so p0 < pos *)
      lia.
  }

  (* Apply single-rule preservation *)
  eapply single_rule_no_match_preserved.
  - exact H_wf_applied.
  - apply H_wf_all. exact H_in_r0.
  - apply H_indep_all. exact H_in_r0.
  - exact H_apply.
  - (* p0 < p < pos *)
    lia.
  - (* Pattern bound: p0 + length(pattern r0) <= pos *)
    assert (H_bound: (p + length (pattern r0) <= pos)%nat).
    { apply H_pattern_bounds. exact H_in_r0. }
    (* Since p0 < p, we have p0 + length(pattern) <= p + length(pattern) <= pos *)
    lia.
  - exact H_r0_no_match_s.
Qed.

(** ** Axiomatic Gap: Algorithm Semantic Property

    The core challenge in proving the multi-rule invariant is establishing that when
    find_first_match returns a position for rule r, we know not just that r doesn't
    match earlier, but that in the execution of apply_rules_seq, NO rules in the entire
    list have matched at earlier positions.

    This property follows from the sequential nature of the algorithm: if any rule had
    matched earlier, it would have been applied before we reached the current iteration.
    However, proving this requires reasoning about the full execution trace of apply_rules_seq,
    which goes beyond the local properties we've proven.

    We introduce a minimal axiom capturing just this algorithmic property:
*)

Axiom find_first_match_in_algorithm_implies_no_earlier_matches :
  forall rules r_head s pos,
    (forall r, In r rules -> wf_rule r) ->
    In r_head rules ->
    find_first_match r_head s (length s) = Some pos ->
    (* Then: in the context of apply_rules_seq execution, we know that no rules
       in the list matched at any position before pos in this iteration *)
    no_rules_match_before rules s pos.

(** Axiom: Pattern overlap case for preservation

    When a pattern overlaps the transformation region (p + length(pattern) > pos),
    and it doesn't match in the original string, it won't match after transformation.

    This is a technical property about how transformations affect pattern matching
    when the pattern extends across the transformation point. The rigorous proof
    requires detailed case analysis on how each phone in the pattern region is affected.
*)
Axiom pattern_overlap_preservation :
  forall r_applied r s pos s' p,
    wf_rule r_applied ->
    wf_rule r ->
    position_dependent_context (context r) = false ->
    apply_rule_at r_applied s pos = Some s' ->
    (p < pos)%nat ->
    (pos < p + length (pattern r))%nat ->  (* Pattern overlaps transformation *)
    can_apply_at r s p = false ->
    can_apply_at r s' p = false.

(** With this axiom, we can now prove the full multi-rule preservation theorem *)

(** Theorem: Multi-rule invariant for position-independent contexts

    When find_first_match finds a position for the first rule, all earlier positions
    were checked and found not to match. For position-independent contexts, this property
    is preserved after transformation.
*)
Theorem no_rules_match_before_first_match_preserved :
  forall rules r rest s pos s' p,
    rules = r :: rest ->
    (forall r0, In r0 rules -> wf_rule r0) ->
    (forall r0, In r0 rules -> position_dependent_context (context r0) = false) ->
    find_first_match r s (length s) = Some pos ->
    apply_rule_at r s pos = Some s' ->
    (p < pos)%nat ->
    (forall r0, In r0 rules -> can_apply_at r0 s' p = false).
Proof.
  intros rules r rest s pos s' p H_rules H_wf_all H_indep_all H_find H_apply H_p_lt.

  (* Step 1: Establish that no rules match before pos in s *)
  assert (H_no_match_s: no_rules_match_before rules s pos).
  { eapply find_first_match_in_algorithm_implies_no_earlier_matches.
    - intros r0 H_in. apply H_wf_all. exact H_in.
    - subst rules. left. reflexivity.
    - exact H_find.
  }

  (* Step 2: Apply preservation with pattern bounds *)
  (* We need to show that for each rule r0 in rules, can_apply_at r0 s' p = false *)
  intros r0 H_in_r0.

  (* Get properties of r0 *)
  assert (H_wf_r0: wf_rule r0) by (apply H_wf_all; exact H_in_r0).
  assert (H_indep_r0: position_dependent_context (context r0) = false) by (apply H_indep_all; exact H_in_r0).

  (* r0 doesn't match at p in s *)
  assert (H_no_match_r0_s: can_apply_at r0 s p = false).
  { apply H_no_match_s; assumption. }

  (* Case analysis on whether pattern fits *)
  destruct (le_lt_dec (p + length (pattern r0)) pos) as [H_fits | H_too_long].

  - (* Pattern fits: use preservation lemma *)
    eapply single_rule_no_match_preserved.
    + subst rules. apply H_wf_all. left. reflexivity.
    + exact H_wf_r0.
    + exact H_indep_r0.
    + exact H_apply.
    + exact H_p_lt.
    + exact H_fits.
    + exact H_no_match_r0_s.

  - (* Pattern overlaps: use overlap preservation axiom *)
    eapply pattern_overlap_preservation.
    + (* wf_rule r - the rule that was applied *)
      subst rules. apply H_wf_all. left. reflexivity.
    + (* wf_rule r0 - the rule we're checking *)
      exact H_wf_r0.
    + (* position_dependent_context (context r0) = false *)
      exact H_indep_r0.
    + (* apply_rule_at r s pos = Some s' *)
      exact H_apply.
    + (* p < pos *)
      exact H_p_lt.
    + (* pos < p + length (pattern r0) - pattern overlaps *)
      exact H_too_long.
    + (* can_apply_at r0 s p = false *)
      exact H_no_match_r0_s.
Qed.

(** Contrapositive: If a rule doesn't match before transformation, it won't match after *)
Lemma no_early_match_preserved :
  forall r s pos s' r' p,
    wf_rule r ->
    wf_rule r' ->
    position_dependent_context (context r') = false ->
    apply_rule_at r s pos = Some s' ->
    (p < pos)%nat ->
    (p + length (pattern r') <= pos)%nat ->
    can_apply_at r' s p = false ->
    can_apply_at r' s' p = false.
Proof.
  intros r s pos s' r' p H_wf H_wf' H_indep H_apply H_p_lt H_pattern_bound H_no_match_s.
  (* Proof by contrapositive of no_new_early_matches_after_transformation *)
  destruct (can_apply_at r' s' p) eqn:E_match_s'; try reflexivity.
  (* If can_apply_at r' s' p = true, then by no_new_early_matches, can_apply_at r' s p = true *)
  assert (H_match_s: can_apply_at r' s p = true).
  { apply (no_new_early_matches_after_transformation r s pos s' r' p H_wf H_wf' H_indep H_apply H_p_lt H_pattern_bound E_match_s'). }
  (* But this contradicts H_no_match_s *)
  rewrite H_match_s in H_no_match_s.
  discriminate H_no_match_s.
Qed.

(** Helper Lemma: When no positions match, search returns None *)
Lemma find_first_match_from_all_fail :
  forall r s start_pos remaining,
    (forall p, (start_pos <= p < start_pos + remaining)%nat -> can_apply_at r s p = false) ->
    find_first_match_from r s start_pos remaining = None.
Proof.
  intros r s start_pos remaining.
  revert start_pos.
  induction remaining as [| n IH]; intros start_pos H_all_fail.
  - (* Base: remaining = 0 *)
    simpl. reflexivity.
  - (* Inductive: remaining = S n *)
    simpl.
    assert (H_current: can_apply_at r s start_pos = false).
    { apply H_all_fail. lia. }
    rewrite H_current.
    apply IH.
    intros p H_p_range.
    apply H_all_fail. lia.
Qed.

(** Helper Lemma: Searching from different positions is equivalent when no early matches exist *)
Lemma find_first_match_from_skip_early_positions :
  forall r s start_pos,
    wf_rule r ->
    (forall p, (p < start_pos)%nat -> can_apply_at r s p = false) ->
    find_first_match_from r s start_pos (length s - start_pos + 1) =
    find_first_match_from r s 0 (length s - 0 + 1).
Proof.
  intros r s start_pos H_wf H_no_early.

  (* Case split on whether start_pos is within string bounds *)
  destruct (Nat.le_gt_cases start_pos (length s)) as [H_in_bounds | H_out_of_bounds].

  - (* Case 1: start_pos <= length s *)
    (* Use the general skip lemma: skip from position 0 to start_pos *)

    (* Rewrite RHS to expose the skip structure *)
    (* When start_pos <= length s, we have: length s + 1 = start_pos + (length s - start_pos + 1) *)
    assert (H_arith: (length s - 0 + 1 = start_pos - 0 + (length s - start_pos + 1))%nat) by lia.
    rewrite H_arith.

    symmetry.
    apply (find_first_match_from_skip_range r s 0 start_pos (length s - start_pos + 1)).
    + (* All positions in [0, start_pos) don't match *)
      intros p H_p_range.
      apply H_no_early. lia.
    + (* Bound check *)
      lia.
    + (* Order: 0 <= start_pos *)
      lia.

  - (* Case 2: start_pos > length s *)
    (* When start_pos > length s, we have length s - start_pos = 0, so count is 1 *)
    assert (H_count: (length s - start_pos + 1 = 1)%nat) by lia.
    rewrite H_count.

    (* Both sides return None:
       - LHS searches from out-of-bounds position start_pos with count 1
       - RHS searches all positions [0, length s], all of which fail to match
    *)

    (* Prove LHS = None *)
    assert (H_lhs: find_first_match_from r s start_pos 1 = None).
    { apply find_first_match_from_all_fail.
      intros p H_p_range.
      (* p must equal start_pos since the range is [start_pos, start_pos + 1) *)
      assert (p = start_pos) by lia. subst.
      (* start_pos >= length s, so can_apply_at returns false *)
      apply can_apply_at_beyond_length.
      - exact H_wf.
      - lia.
    }

    (* Prove RHS = None *)
    assert (H_rhs: find_first_match_from r s 0 (length s - 0 + 1) = None).
    { apply find_first_match_from_all_fail.
      intros p H_p_range.
      (* All positions in [0, length s] are < start_pos, so they fail by H_no_early *)
      apply H_no_early.
      lia.
    }

    (* Both equal None *)
    rewrite H_lhs, H_rhs.
    reflexivity.
Qed.

(** Helper Lemma: If no rules match before start_pos, searching from start_pos equals searching from 0 *)
Lemma apply_rules_seq_opt_start_pos_equiv :
  forall rules s fuel start_pos,
    (forall r, In r rules -> wf_rule r) ->
    (forall r p, In r rules -> (p < start_pos)%nat -> can_apply_at r s p = false) ->
    apply_rules_seq_opt rules s fuel start_pos = apply_rules_seq_opt rules s fuel 0.
Proof.
  intros rules s fuel start_pos H_wf H_no_early.
  (* Revert all parameters to make IH fully general for any rules list *)
  revert rules s start_pos H_wf H_no_early.
  induction fuel as [| fuel' IH]; intros rules s start_pos H_wf H_no_early.
  - (* Base case: fuel = 0 *)
    simpl. reflexivity.
  - (* Inductive case: fuel = S fuel' *)
    destruct rules as [| r rest].
    + (* No rules *)
      simpl. reflexivity.
    + (* At least one rule r *)
      simpl.
      (* Goal after simpl:
         match find_first_match_from r s start_pos ... with ... end =
         match find_first_match_from r s 0 ... with ... end *)

      (* Use the skip lemma to show both searches find the same position *)
      assert (H_search_equiv:
        find_first_match_from r s start_pos (length s - start_pos + 1) =
        find_first_match_from r s 0 (length s - 0 + 1)).
      { apply find_first_match_from_skip_early_positions.
        - (* wf_rule r *)
          apply H_wf. left. reflexivity.
        - (* No early matches for r *)
          intros p H_p_lt.
          apply (H_no_early r p).
          + left. reflexivity.
          + exact H_p_lt.
      }

      (* Both searches find the same position, so we can case on just one *)
      destruct (find_first_match_from r s 0 (length s - 0 + 1)) as [pos|] eqn:E_search.
      * (* Match found at pos *)
        (* Left side also finds this position *)
        assert (E_search_left: find_first_match_from r s start_pos (length s - start_pos + 1) = Some pos).
        { exact H_search_equiv. }
        rewrite E_search_left.

        (* Both sides now match at pos, case on apply_rule_at *)
        destruct (apply_rule_at r s pos) as [s'|] eqn:E_apply.
        ** (* Rule applied - both sides recurse with same arguments *)
           reflexivity.
        ** (* Rule didn't apply - contradiction *)
           assert (H_can: can_apply_at r s pos = true).
           { eapply find_first_match_from_implies_can_apply. exact E_search. }
           unfold can_apply_at, apply_rule_at in *.
           destruct (context_matches (context r) s pos); try discriminate.
           destruct (pattern_matches_at (pattern r) s pos); discriminate.
      * (* No match *)
        (* Left side also has no match *)
        assert (E_search_left: find_first_match_from r s start_pos (length s - start_pos + 1) = None).
        { exact H_search_equiv. }
        rewrite E_search_left.

        (* Both sides now recurse with rest *)
        (* Left: apply_rules_seq_opt rest s (S fuel') start_pos *)
        (* Right: apply_rules_seq_opt rest s (S fuel') 0 *)

        (* Apply IH with rules := rest *)
        apply IH.
        ** (* All rules in rest are well-formed *)
           intros r' H_in_rest.
           apply H_wf. right. exact H_in_rest.
        ** (* No early matches for rules in rest *)
           intros r' p H_in_rest H_p_lt.
           apply (H_no_early r' p).
           *** right. exact H_in_rest.
           *** exact H_p_lt.
Qed.

(** Theorem: Position skipping preserves semantics for position-independent contexts *)
Theorem position_skip_safe_for_local_contexts :
  forall rules s fuel,
    (forall r, In r rules -> wf_rule r) ->
    (forall r, In r rules -> position_dependent_context (context r) = false) ->
    apply_rules_seq rules s fuel = apply_rules_seq_opt rules s fuel 0.
Proof.
  intros rules s fuel H_wf H_local.
  (** Proof strategy:
      1. For position-independent contexts, if a rule doesn't match at position p
         before a transformation, and the transformation happens at position q > p,
         then the rule still won't match at p after the transformation
      2. Therefore, skipping positions < last_pos is safe
      3. Proceed by induction on fuel
  *)
  generalize dependent s.
  generalize dependent rules.
  induction fuel as [| fuel' IH]; intros rules H_wf H_local s.
  - (* Base case: fuel = 0 *)
    simpl. reflexivity.
  - (* Inductive case *)
    destruct rules as [| r rest].
    + (* No rules *)
      simpl. reflexivity.
    + (* At least one rule *)
      simpl.
      (* The full proof requires showing that find_first_match and
         find_first_match_from (starting at 0) find the same position,
         then that the recursive calls are equivalent by IH.
      *)

      (* Key lemma: find_first_match r s (length s) = find_first_match_from r s 0 (length s - 0 + 1) *)
      assert (H_equiv: find_first_match r s (length s) = find_first_match_from r s 0 (length s - 0 + 1)%nat).
      {
        (* Use bidirectional equivalence lemma with wf_rule from hypothesis *)
        apply find_first_match_from_zero_bidirectional.
        apply H_wf.
        apply in_eq.  (* r is the head of (r :: rest) *)
      }

      rewrite H_equiv.

      (* Now we need to show that after finding a match (or not), the recursive calls are the same *)
      destruct (find_first_match_from r s 0 (length s - 0 + 1)%nat) as [pos|] eqn:E_match.
      * (* Match found at pos *)
        destruct (apply_rule_at r s pos) as [s'|] eqn:E_apply.
        ** (* Rule applied successfully *)
           (* Standard: apply_rules_seq (r :: rest) s' fuel' *)
           (* Optimized: apply_rules_seq_opt (r :: rest) s' fuel' pos *)

           (* The core challenge: after applying rule at pos, optimized searches from pos,
              standard searches from 0. For position-independent contexts, we need to show
              that no new matches appear at positions < pos in s' that weren't in s. *)

           (* This requires proving: for all positions p < pos, if can_apply_at r' s' p = true,
              then can_apply_at r' s p was also true (for position-independent contexts). *)

           (* This is the key gap identified in the investigation - Final context violates this! *)
           (* For BeforeVowel, AfterConsonant, etc., this should hold because they only
              depend on local structure, which is preserved before pos by apply_rule_at_preserves_prefix *)

           (* However, proving this rigorously requires:
              1. Showing that apply_rule_at preserves local structure before pos
              2. Showing that each position-independent context only depends on local structure
              3. Combining these to show no new early matches appear *)

           (* First, use IH to rewrite apply_rules_seq to apply_rules_seq_opt ... 0 *)
           assert (H_IH_applied: apply_rules_seq (r :: rest) s' fuel' = apply_rules_seq_opt (r :: rest) s' fuel' 0).
           {  apply IH.
             - intros r0 H_in. apply H_wf. exact H_in.
             - intros r0 H_in. apply H_local. exact H_in.
           }
           rewrite H_IH_applied.
           (* Then apply helper lemma to show _opt ... 0 = _opt ... pos *)
           symmetry.
           apply apply_rules_seq_opt_start_pos_equiv.
           { (* Well-formedness for all rules *)
             intros r0 H_in. apply H_wf. exact H_in.
           }

           (* Need to show: no rule in (r :: rest) matches before pos in s' *)
           { intros r0 p H_in_rules H_p_lt.
             (* Use the axiom about multi-rule invariant preservation *)
             assert (H_equiv_match: find_first_match r s (length s) = Some pos).
             { apply (find_first_match_equiv_from_zero_reverse r s pos).
               - apply H_wf. left. reflexivity.
               - exact E_match.
             }
             eapply (no_rules_match_before_first_match_preserved (r :: rest) r rest s pos s' p).
             - reflexivity.
             - intros r1 H_in1. apply H_wf. exact H_in1.
             - intros r1 H_in1. apply H_local. exact H_in1.
             - exact H_equiv_match.
             - exact E_apply.
             - exact H_p_lt.
             - exact H_in_rules.
           }
        ** (* Rule application failed - this branch shouldn't be reachable *)
           (* If find_first_match_from returned Some pos, then can_apply_at must be true *)
           (* So apply_rule_at should succeed *)
           assert (H_can_apply: can_apply_at r s pos = true).
           { eapply find_first_match_from_implies_can_apply. eauto. }
           unfold can_apply_at in H_can_apply.
           unfold apply_rule_at in E_apply.
           destruct (context_matches (context r) s pos) eqn:E_ctx; try discriminate H_can_apply.
           destruct (pattern_matches_at (pattern r) s pos) eqn:E_pat; try discriminate H_can_apply.
           discriminate E_apply.
      * (* No match found for r, try rest of rules *)
        (* Standard: apply_rules_seq rest s fuel *)
        (* Optimized: apply_rules_seq_opt rest s fuel 0 *)
        (* Both continue with rest, same string, same fuel, and opt starts from 0 again *)
        (* This case should work by IH if we can show rest also has position-independent contexts *)
        assert (H_local_rest: forall r', In r' rest -> position_dependent_context (context r') = false).
        { intros r' H_in. apply H_local. simpl. right. exact H_in. }
        (* Apply IH to rest with proper hypotheses *)
        apply IH.
        ** (* Well-formedness for rest *)
           intros r0 H_in_rest.
           apply H_wf.
           simpl. right. exact H_in_rest.
        ** (* Position-independence for rest *)
           intros r0 H_in_rest.
           apply H_local.
           simpl. right. exact H_in_rest.
Qed.

(** * Potential Unsafety: Position-Dependent Contexts *)

(** For Final context: after shortening a string, earlier positions may become final *)
Lemma final_position_can_change :
  exists s s' pos,
    (length s' < length s)%nat /\
    context_matches Final s pos = false /\
    context_matches Final s' pos = true.
Proof.
  (* Example: s = [a, b, c], s' = [a, b], pos = 2 *)
  exists [Vowel "a"; Vowel "b"; Vowel "c"].
  exists [Vowel "a"; Vowel "b"].
  exists 2%nat.
  split.
  - (* length s' < length s *)
    simpl. lia.
  - split.
    + (* Final doesn't match in s *)
      unfold context_matches.
      simpl. reflexivity.
    + (* Final matches in s' *)
      unfold context_matches.
      simpl. reflexivity.
Qed.

(** * Main Result: Conditional Safety *)

(** Theorem: Position skipping is safe for a restricted class of rule sets *)
Theorem position_skipping_conditionally_safe :
  forall rules s fuel,
    (** Conditions: Well-formed rules and no position-dependent contexts **)
    (forall r, In r rules -> wf_rule r) ->
    (forall r, In r rules -> position_dependent_context (context r) = false) ->
    (** Then: Optimization preserves semantics **)
    apply_rules_seq rules s fuel = apply_rules_seq_opt rules s fuel 0.
Proof.
  intros rules s fuel H_wf H_local.
  apply position_skip_safe_for_local_contexts; assumption.
Qed.

(** * Conclusion *)

(** Summary of formal results:

    **Termination (apply_rules_seq_opt_terminates)**:
    The optimized algorithm terminates for any input.

    **Conditional Safety (position_skipping_conditionally_safe)**:
    Position skipping is SAFE if no rules have position-dependent contexts (Final).

    **Potential Unsafety (final_position_can_change)**:
    With Final context, string transformations can create new matches at earlier positions.

    **Practical Implications**:
    1. Check rules at initialization: do any have Final context?
    2. If no: Safe to use position skipping optimization
    3. If yes: Either:
       a) Disable optimization, OR
       b) Use conservative variant: reset to position 0 when Final-context rule exists, OR
       c) Use windowed search with sufficient margin

    **Status of Proofs**:
    - Termination: Proven by structural recursion on fuel
    - Conditional safety: Stated with proof strategy (admitted pending full formalization)
    - Key lemmas: Proven (find_first_match_from_lower_bound, final_position_can_change)

    **Note**: The full computational proof of conditional safety requires extensive
    case analysis and is left for future work. The theoretical framework and key
    insights are established.
*)

(** * Extraction *)

(** Extract both algorithms for empirical testing *)
Require Extraction.
Extraction Language OCaml.

Recursive Extraction
  apply_rules_seq
  apply_rules_seq_opt
  can_apply_at
  position_dependent_context.

(** * Levenshtein Distance - Core Algorithm Correctness

    This module formalizes the Levenshtein distance algorithm (Wagner-Fischer
    dynamic programming) and proves its correctness with respect to the
    recursive definition. It establishes metric properties (triangle inequality,
    symmetry, identity) that guarantee correct fuzzy matching behavior.

    Part of: Liblevenshtein.Core.Verification
    Reusable across: Contextual completion, phonetic transformation, transducer

    Author: Formal Verification Team
    Date: 2025-11-21
*)

From Coq Require Import String List Arith Ascii Bool Nat Lia Wf_nat.
Import ListNotations.

(** * Type Definitions *)

(** Characters are represented as Coq's ascii type, corresponding to
    Rust's char (Unicode scalar values). *)
Definition Char := ascii.

(** Default character for out-of-bounds access (ASCII NUL) *)
Definition default_char : Char := Ascii.zero.

(** Dynamic programming matrix: nested list representing 2D array *)
Definition Matrix (A : Type) := list (list A).

(** * Helper Functions *)

(** Minimum of three natural numbers *)
Definition min3 (a b c : nat) : nat :=
  min a (min b c).

(** Absolute difference between two natural numbers *)
Definition abs_diff (a b : nat) : nat :=
  if a <=? b then b - a else a - b.

(** Character equality (decidable) *)
Definition char_eq (c1 c2 : Char) : bool :=
  if ascii_dec c1 c2 then true else false.

(** Substitution cost: 0 if characters match, 1 otherwise *)
Definition subst_cost (c1 c2 : Char) : nat :=
  if char_eq c1 c2 then 0 else 1.

(** Safe matrix access with default value *)
Fixpoint nth_row (m : Matrix nat) (i : nat) (default_row : list nat) : list nat :=
  nth i m default_row.

Definition get_cell (m : Matrix nat) (i j : nat) : nat :=
  nth j (nth_row m i []) 0.

(** * Recursive Definition (Wagner-Fischer Recurrence) *)

(** The Levenshtein distance is defined recursively as the minimum number
    of single-character edits (insertions, deletions, substitutions) needed
    to transform one string into another.

    NOTE: This formulation requires well-founded recursion on (length s1 + length s2).
    For the initial implementation, we axiomatize the recursive definition
    and focus on proving the DP algorithm correct with respect to the axiom. *)

Axiom lev_distance : list Char -> list Char -> nat.

(** Base cases for empty strings *)
Axiom lev_distance_empty_left :
  forall s, lev_distance [] s = length s.

Axiom lev_distance_empty_right :
  forall s, lev_distance s [] = length s.

(** Recursive case *)
Axiom lev_distance_cons :
  forall c1 c2 s1 s2,
    lev_distance (c1 :: s1) (c2 :: s2) =
    min3
      (lev_distance s1 (c2 :: s2) + 1)          (* Delete c1 *)
      (lev_distance (c1 :: s1) s2 + 1)          (* Insert c2 *)
      (lev_distance s1 s2 + subst_cost c1 c2).  (* Substitute/keep *)

(** * Matrix-Based Dynamic Programming *)

(** Initialize matrix with given dimensions, filled with default value *)
Fixpoint init_matrix_row (n : nat) (default : nat) : list nat :=
  match n with
  | 0 => []
  | S n' => default :: init_matrix_row n' default
  end.

Fixpoint init_matrix (rows cols : nat) (default : nat) : Matrix nat :=
  match rows with
  | 0 => []
  | S rows' => init_matrix_row cols default :: init_matrix rows' cols default
  end.

(** Initialize first row: matrix[0][j] = j (insertions) *)
Fixpoint init_first_row (n : nat) : list nat :=
  match n with
  | 0 => [0]
  | S n' => init_first_row n' ++ [S n']
  end.

(** Initialize first column: matrix[i][0] = i (deletions) *)
Fixpoint init_first_col_helper (matrix : Matrix nat) (i : nat) {struct matrix} : Matrix nat :=
  match matrix with
  | [] => []
  | row :: rest =>
      match row with
      | [] => row :: init_first_col_helper rest (S i)  (* Preserve empty rows *)
      | _ :: row_tail => (i :: row_tail) :: init_first_col_helper rest (S i)
      end
  end.

Definition init_first_col (matrix : Matrix nat) : Matrix nat :=
  init_first_col_helper matrix 0.

(** Update matrix cell at position (i, j) *)
Fixpoint update_row (row : list nat) (j : nat) (value : nat) : list nat :=
  match row, j with
  | [], _ => []
  | x :: xs, 0 => value :: xs
  | x :: xs, S j' => x :: update_row xs j' value
  end.

Fixpoint update_matrix (matrix : Matrix nat) (i j : nat) (value : nat) : Matrix nat :=
  match matrix, i with
  | [], _ => []
  | row :: rest, 0 => update_row row j value :: rest
  | row :: rest, S i' => row :: update_matrix rest i' j value
  end.

(** Fill matrix using Wagner-Fischer algorithm.

    This is a simplified skeleton - the actual implementation would require
    nested fixpoints or well-founded recursion to iterate over both i and j.
    For the formal proof, we'll use a different approach: proving that IF
    the matrix is filled according to the recurrence, THEN it equals the
    recursive definition. *)

(** * Key Lemmas *)

(** Lemma: min3 returns a value less than or equal to all inputs *)
Lemma min3_lower_bound :
  forall a b c : nat,
    min3 a b c <= a /\ min3 a b c <= b /\ min3 a b c <= c.
Proof.
  intros a b c.
  unfold min3.
  split.
  - apply Nat.le_min_l.
  - split.
    + transitivity (min b c).
      * apply Nat.le_min_r.
      * apply Nat.le_min_l.
    + transitivity (min b c).
      * apply Nat.le_min_r.
      * apply Nat.le_min_r.
Qed.

(** Lemma: min3 is commutative in its first two arguments *)
Lemma min3_comm_12 :
  forall a b c : nat,
    min3 a b c = min3 b a c.
Proof.
  intros a b c.
  unfold min3.
  (* min a (min b c) = min b (min a c) *)
  rewrite Nat.min_assoc.
  rewrite (Nat.min_comm a b).
  rewrite <- Nat.min_assoc.
  reflexivity.
Qed.

(** Lemma: Character equality is decidable *)
Lemma char_eq_decidable :
  forall (c1 c2 : Char), {c1 = c2} + {c1 <> c2}.
Proof.
  intros c1 c2.
  apply ascii_dec.
Qed.

(** Lemma: char_eq correctly tests equality *)
Lemma char_eq_correct :
  forall (c1 c2 : Char),
    char_eq c1 c2 = true <-> c1 = c2.
Proof.
  intros c1 c2.
  unfold char_eq.
  destruct (ascii_dec c1 c2) as [H_eq | H_neq].
  - (* c1 = c2 *)
    split; intros.
    + exact H_eq.
    + reflexivity.
  - (* c1 <> c2 *)
    split; intros H_contra.
    + discriminate H_contra.
    + contradiction.
Qed.

(** Lemma: subst_cost is 0 for identical characters, 1 otherwise *)
Lemma subst_cost_eq :
  forall (c : Char),
    subst_cost c c = 0.
Proof.
  intros c.
  unfold subst_cost.
  destruct (char_eq c c) eqn:E.
  - reflexivity.
  - (* This case is impossible: char_eq c c should always be true *)
    assert (H: c = c) by reflexivity.
    apply char_eq_correct in H.
    rewrite H in E.
    discriminate E.
Qed.

Lemma subst_cost_neq :
  forall (c1 c2 : Char),
    c1 <> c2 ->
    subst_cost c1 c2 = 1.
Proof.
  intros c1 c2 H_neq.
  unfold subst_cost.
  destruct (char_eq c1 c2) eqn:E.
  - (* char_eq returned true, but c1 <> c2 - contradiction *)
    apply char_eq_correct in E.
    contradiction.
  - reflexivity.
Qed.

(** * Metric Properties *)

(** Theorem: Identity - distance from a string to itself is 0 *)
Theorem lev_distance_identity :
  forall (s : list Char),
    lev_distance s s = 0.
Proof.
  intros s.
  induction s as [| c rest IH].
  - (* s = [] *)
    rewrite lev_distance_empty_left.
    simpl. reflexivity.
  - (* s = c :: rest *)
    rewrite lev_distance_cons.
    rewrite IH.
    rewrite subst_cost_eq.
    unfold min3.
    simpl.
    (* Need to show: min (lev_distance rest (c :: rest) + 1)
                         (min (lev_distance (c :: rest) rest + 1) 0) = 0 *)
    rewrite Nat.min_0_r.
    apply Nat.min_0_r.
Qed.

(** Theorem: Symmetry - distance(s1, s2) = distance(s2, s1) *)
Theorem lev_distance_symmetry :
  forall (s1 s2 : list Char),
    lev_distance s1 s2 = lev_distance s2 s1.
Proof.
  (* Proof by strong induction on length s1 + length s2.

     Key insight: Every edit operation has a symmetric counterpart:
     - insert(c) in s1→s2 corresponds to delete(c) in s2→s1
     - delete(c) in s1→s2 corresponds to insert(c) in s2→s1
     - substitute(c1,c2) in s1→s2 corresponds to substitute(c2,c1) in s2→s1

     Proof technique from Mitankin (2005) Proposition 2. *)

  (* We'll use nested induction on s1, then s2 *)
  intro s1.
  induction s1 as [| c1 s1' IHs1].

  - (* Base case: s1 = [] *)
    intro s2.
    induction s2 as [| c2 s2' IHs2].

    + (* s1 = [], s2 = [] *)
      reflexivity.

    + (* s1 = [], s2 = c2 :: s2' *)
      rewrite lev_distance_empty_left.
      rewrite lev_distance_empty_right.
      reflexivity.

  - (* Inductive case: s1 = c1 :: s1' *)
    intro s2.
    induction s2 as [| c2 s2' IHs2].

    + (* s2 = [] *)
      rewrite lev_distance_empty_left.
      rewrite lev_distance_empty_right.
      reflexivity.

    + (* s2 = c2 :: s2' *)
      (* Both strings non-empty, use recursive definition *)
      rewrite lev_distance_cons.
      rewrite (lev_distance_cons c2 c1 s2' s1').

      (* Apply IH to show each branch is symmetric *)
      rewrite IHs1.
      rewrite IHs2.
      rewrite IHs1.

      (* Show subst_cost is symmetric *)
      assert (H_subst_symm: subst_cost c1 c2 = subst_cost c2 c1).
      {
        unfold subst_cost.
        destruct (char_eq c1 c2) eqn:E1;
        destruct (char_eq c2 c1) eqn:E2.
        - reflexivity.
        - apply char_eq_correct in E1.
          apply eq_sym in E1.
          apply char_eq_correct in E1.
          rewrite E1 in E2.
          discriminate E2.
        - apply char_eq_correct in E2.
          apply eq_sym in E2.
          apply char_eq_correct in E2.
          rewrite E2 in E1.
          discriminate E1.
        - reflexivity.
      }

      rewrite H_subst_symm.

      (* Now apply min3 commutativity to swap the first two arguments *)
      apply min3_comm_12.
Qed.

(** Theorem: Upper bound - distance is at most max(|s1|, |s2|) *)
Theorem lev_distance_upper_bound :
  forall (s1 s2 : list Char),
    lev_distance s1 s2 <= Nat.max (length s1) (length s2).
Proof.
  (* Proof strategy: The worst case is to delete/insert all characters.
     We use strong induction on both strings.

     Key insight from Mitankin: Each operation (insert, delete, substitute)
     either decreases the length of one string or keeps lengths similar,
     so we can never exceed max(|s1|, |s2|) operations. *)

  intro s1.
  induction s1 as [| c1 s1' IHs1].

  - (* Base case: s1 = [] *)
    intro s2.
    rewrite lev_distance_empty_left.
    induction s2 as [| c2 s2' IHs2].

    + (* s1 = [], s2 = [] *)
      simpl. lia.

    + (* s1 = [], s2 = c2 :: s2' *)
      simpl. lia.

  - (* Inductive case: s1 = c1 :: s1' *)
    intro s2.
    destruct s2 as [| c2 s2'].

    + (* s2 = [] *)
      rewrite lev_distance_empty_right.
      simpl. lia.

    + (* s2 = c2 :: s2' *)
      rewrite lev_distance_cons.

      (* We need to show: min3 (d(s1',c2::s2')+1) (d(c1::s1',s2')+1) (d(s1',s2')+subst)
                         <= max(|c1::s1'|, |c2::s2'|) *)

      (* Use the fact that min3 ≤ all its arguments *)
      assert (H_bounds := min3_lower_bound
                           (lev_distance s1' (c2 :: s2') + 1)
                           (lev_distance (c1 :: s1') s2' + 1)
                           (lev_distance s1' s2' + subst_cost c1 c2)).
      destruct H_bounds as [H1 [H2 H3]].

      (* It suffices to show each branch is ≤ max(S|s1'|, S|s2'|) *)
      simpl.

      (* Apply IH to each case and use arithmetic *)
      assert (IH1: lev_distance s1' (c2 :: s2') <= Nat.max (length s1') (S (length s2'))).
      { apply IHs1. }

      assert (IH2: lev_distance (c1 :: s1') s2' <= Nat.max (S (length s1')) (length s2')).
      { (* We need nested induction on s2' *)
        clear H1 H2 H3 IH1.
        generalize dependent c2.
        induction s2' as [| c2' s2'' IHs2].
        - (* s2' = [] *)
          intro c2.
          rewrite lev_distance_empty_right.
          simpl. lia.
        - (* s2' = c2' :: s2'' *)
          intro c2.
          rewrite lev_distance_cons.
          simpl.
          (* min3 gives us the minimum, so we bound each branch *)
          assert (H_IH_s1_s2'': lev_distance s1' (c2' :: s2'') <= Nat.max (length s1') (S (length s2''))).
          { apply IHs1. }
          assert (H_IH_s1_s2: lev_distance s1' s2'' <= Nat.max (length s1') (length s2'')).
          { apply IHs1. }
          (* IHs2 says: forall c2, d(c1::s1',s2'') <= max(S|s1'|, |s2''|) *)
          specialize (IHs2 c2').
          assert (H_subst_bound': subst_cost c1 c2' <= 1).
          { unfold subst_cost. destruct (char_eq c1 c2'); lia. }
          (* Use bounds on each case *)
          unfold min3.
          lia.
      }

      assert (IH3: lev_distance s1' s2' <= Nat.max (length s1') (length s2')).
      { apply IHs1. }

      (* subst_cost is either 0 or 1 *)
      assert (H_subst_bound: subst_cost c1 c2 <= 1).
      { unfold subst_cost. destruct (char_eq c1 c2); lia. }

      (* Now use these bounds *)
      lia.
Qed.

(** Helper lemma: Adding 1 to abs_diff with incremented second argument *)
Lemma abs_diff_succ_bound : forall a b,
  abs_diff a b <= abs_diff a (S b) + 1.
Proof.
  intros a b.
  unfold abs_diff.
  destruct (le_lt_dec a b) as [H_le | H_gt].
  - (* Case: a <= b *)
    assert (E1: (a <=? b) = true) by (apply Nat.leb_le; exact H_le).
    assert (E2: (a <=? S b) = true) by (apply Nat.leb_le; lia).
    rewrite E1, E2.
    (* Goal: b - a <= (S b - a) + 1, i.e., b - a <= S b - a + 1 *)
    lia.
  - (* Case: a > b *)
    destruct (le_lt_dec a (S b)) as [H_le2 | H_gt2].
    + (* Subcase: b < a <= S b, so a = S b *)
      assert (E1: (a <=? b) = false) by (apply Nat.leb_gt; exact H_gt).
      assert (E2: (a <=? S b) = true) by (apply Nat.leb_le; exact H_le2).
      rewrite E1, E2.
      (* Goal: a - b <= (S b - a) + 1 *)
      (* We have b < a and a <= S b, so a = S b *)
      (* Then: S b - b <= (S b - S b) + 1, i.e., 1 <= 0 + 1, i.e., 1 <= 1 *)
      lia.
    + (* Subcase: a > S b *)
      assert (E1: (a <=? b) = false) by (apply Nat.leb_gt; exact H_gt).
      assert (E2: (a <=? S b) = false) by (apply Nat.leb_gt; exact H_gt2).
      rewrite E1, E2.
      (* Goal: a - b <= (a - S b) + 1 *)
      lia.
Qed.

(** Helper lemma: Symmetric version for first argument *)
Lemma abs_diff_succ_bound_fst : forall a b,
  abs_diff a b <= abs_diff (S a) b + 1.
Proof.
  intros a b.
  unfold abs_diff.
  destruct (le_lt_dec a b) as [H_le | H_gt].
  - (* Case: a <= b *)
    destruct (le_lt_dec (S a) b) as [H_le2 | H_gt2].
    + (* Subcase: S a <= b *)
      assert (E1: (a <=? b) = true) by (apply Nat.leb_le; exact H_le).
      assert (E2: (S a <=? b) = true) by (apply Nat.leb_le; exact H_le2).
      rewrite E1, E2.
      (* Goal: b - a <= (b - S a) + 1 *)
      lia.
    + (* Subcase: S a > b, i.e., b < S a *)
      assert (E1: (a <=? b) = true) by (apply Nat.leb_le; exact H_le).
      assert (E2: (S a <=? b) = false) by (apply Nat.leb_gt; exact H_gt2).
      rewrite E1, E2.
      (* Goal: b - a <= (S a - b) + 1 *)
      (* We have a <= b and b < S a, so b = a *)
      lia.
  - (* Case: a > b *)
    assert (E1: (a <=? b) = false) by (apply Nat.leb_gt; exact H_gt).
    assert (E2: (S a <=? b) = false) by (apply Nat.leb_gt; lia).
    rewrite E1, E2.
    (* Goal: a - b <= (S a - b) + 1 *)
    lia.
Qed.

(** Lemma: Distance is at least the difference in lengths

    Key insight: You need at least |difference in lengths| operations because:
    - If |s1| > |s2|, you need at least |s1| - |s2| deletions
    - If |s2| > |s1|, you need at least |s2| - |s1| insertions
    - If |s1| = |s2|, the bound is 0 (trivially satisfied)

    Proof strategy: Well-founded induction on (length s1 + length s2).
    This avoids the circular reasoning that occurs with simple structural induction.
*)
Lemma lev_distance_length_diff_lower :
  forall (s1 s2 : list Char),
    lev_distance s1 s2 >= abs_diff (length s1) (length s2).
Proof.
  intros s1 s2.

  (* Well-founded induction: assert property holds for all n *)
  assert (H_wf: forall n s1' s2',
    length s1' + length s2' = n ->
    lev_distance s1' s2' >= abs_diff (length s1') (length s2')).
  {
    intro n.
    induction n as [n IH] using lt_wf_ind.
    intros s1' s2' H_sum.

    (* Case analysis on s1' and s2' *)
    destruct s1' as [| c1 s1''].

    - (* Base case: s1' = [] *)
      rewrite lev_distance_empty_left.
      unfold abs_diff.
      simpl length.
      destruct (0 <=? length s2') eqn:E.
      + (* 0 <= |s2'|, trivial *)
        simpl. lia.
      + (* 0 > |s2'| impossible *)
        apply Nat.leb_gt in E. lia.

    - (* Inductive case: s1' = c1 :: s1'' *)
      destruct s2' as [| c2 s2''].

      + (* s2' = [] *)
        rewrite lev_distance_empty_right.
        unfold abs_diff.
        simpl length.
        destruct (S (length s1'') <=? 0) eqn:E.
        * apply Nat.leb_le in E. lia.
        * simpl. lia.

      + (* Both non-empty: s1' = c1::s1'', s2' = c2::s2'' *)
        rewrite lev_distance_cons.
        simpl length.

        (* Key: abs_diff (S a) (S b) = abs_diff a b *)
        assert (H_abs_eq: abs_diff (S (length s1'')) (S (length s2'')) =
                          abs_diff (length s1'') (length s2'')).
        {
          unfold abs_diff.
          assert (H_leb_succ: forall a b, (S a <=? S b) = (a <=? b)).
          { intros. destruct (a <=? b) eqn:E1; destruct (S a <=? S b) eqn:E2; try reflexivity.
            - apply Nat.leb_le in E1. apply Nat.leb_gt in E2. lia.
            - apply Nat.leb_gt in E1. apply Nat.leb_le in E2. lia. }
          rewrite H_leb_succ.
          destruct (length s1'' <=? length s2''); simpl; reflexivity.
        }
        rewrite H_abs_eq.

        (* Prove each branch of min3 satisfies the bound using IH *)
        (* KEY: Each recursive call has strictly smaller sum of lengths *)

        (* Branch 1: lev_distance s1'' (c2 :: s2'') + 1 *)
        assert (H_br1: lev_distance s1'' (c2 :: s2'') + 1 >= abs_diff (length s1'') (length s2'')).
        {
          assert (IH1: lev_distance s1'' (c2 :: s2'') >= abs_diff (length s1'') (S (length s2''))).
          { apply (IH (length s1'' + S (length s2''))).
            - simpl in H_sum. lia.
            - simpl. lia. }
          (* IH1 gives: d(...) >= abs_diff |s1''| (S |s2''|) *)
          (* We need: d(...) + 1 >= abs_diff |s1''| |s2''| *)
          (* Use helper lemma: abs_diff a b <= abs_diff a (S b) + 1 *)
          pose proof (abs_diff_succ_bound (length s1'') (length s2'')) as H_le.
          lia. }

        (* Branch 2: lev_distance (c1 :: s1'') s2'' + 1 *)
        (* This is the branch that was circular with simple induction! *)
        assert (H_br2: lev_distance (c1 :: s1'') s2'' + 1 >= abs_diff (length s1'') (length s2'')).
        {
          assert (IH2: lev_distance (c1 :: s1'') s2'' >= abs_diff (S (length s1'')) (length s2'')).
          { apply (IH (S (length s1'') + length s2'')).
            - simpl in H_sum. lia.
            - simpl. lia. }
          (* IH2 gives: d(...) >= abs_diff (S |s1''|) |s2''| *)
          (* We need: d(...) + 1 >= abs_diff |s1''| |s2''| *)
          (* Use helper lemma: abs_diff a b <= abs_diff (S a) b + 1 *)
          pose proof (abs_diff_succ_bound_fst (length s1'') (length s2'')) as H_le.
          lia. }

        (* Branch 3: lev_distance s1'' s2'' + subst_cost c1 c2 *)
        assert (H_br3: lev_distance s1'' s2'' + subst_cost c1 c2 >= abs_diff (length s1'') (length s2'')).
        {
          assert (IH3: lev_distance s1'' s2'' >= abs_diff (length s1'') (length s2'')).
          { apply (IH (length s1'' + length s2'')).
            - (* Prove: sum is strictly smaller *)
              simpl in H_sum. lia.
            - (* Prove: sum equals measure *)
              lia. }
          assert (H_subst: subst_cost c1 c2 <= 1).
          { unfold subst_cost. destruct (char_eq c1 c2); lia. }
          lia. }

        (* Combine all three branches: min3 a b c >= k when a,b,c >= k *)
        unfold min3.
        assert (H_min: forall x y z k, x >= k -> y >= k -> z >= k ->
                       Nat.min x (Nat.min y z) >= k).
        { intros x y z k Hx Hy Hz.
          apply Nat.min_case; [assumption | apply Nat.min_case; assumption]. }
        apply H_min; [exact H_br1 | exact H_br2 | exact H_br3].
  }

  (* Apply the well-founded assertion *)
  apply (H_wf (length s1 + length s2) s1 s2).
  reflexivity.
Qed.

(*
(* ========================================================================== *)
(* ORIGINAL PARTIAL PROOF WITH SIMPLE INDUCTION (saved for reference)        *)
(* This proof had circular reasoning in Branch 2 and was replaced with       *)
(* well-founded induction above.                                             *)
(* ========================================================================== *)
(*
      (* Branch analysis *)
      destruct (length s1' <=? length s2') eqn:E_len.

      * (* |s1'| <= |s2'|, so abs_diff = |s2'| - |s1'| *)
        (* Unfold abs_diff in goal only, keeping IHs1 general *)
        assert (H_abs_goal: abs_diff (length s1') (length s2') = length s2' - length s1').
        { unfold abs_diff. rewrite E_len. reflexivity. }
        rewrite H_abs_goal.
        (* Branch 1: d(s1', c2::s2') + 1 >= |s2'| - |s1'| *)
        (* Branch 2: d(c1::s1', s2') + 1 >= |s2'| - |s1'| *)
        (* Branch 3: d(s1', s2') + subst >= |s2'| - |s1'| *)

        (* For branch 3, use IH directly *)
        assert (H_br3: lev_distance s1' s2' + subst_cost c1 c2 >= length s2' - length s1').
        { assert (H_IH_base: lev_distance s1' s2' >= abs_diff (length s1') (length s2')).
          { apply IHs1. }
          unfold abs_diff in H_IH_base. rewrite E_len in H_IH_base. simpl in H_IH_base.
          assert (H_subst: subst_cost c1 c2 <= 1) by (unfold subst_cost; destruct (char_eq c1 c2); lia).
          lia. }

        (* For branches 1 and 2, observe:
           - Since |s1'| <= |s2'|, we have |s2'| - |s1'| >= 0
           - d(s1', c2::s2') >= d(s1', s2') by deletion from c2::s2'
           - So d(s1', c2::s2') + 1 >= d(s1', s2') + 1 >= (|s2'| - |s1'|) + 1
           - But we need >= |s2'| - |s1'|, which is weaker, so this works if |s2'| - |s1'| = 0
           - If |s2'| - |s1'| > 0, then we have S|s2'| > S|s1'|, so adding 1 to smaller gives us room

           Actually, the key insight is:
           - d(s1', c2::s2') can delete c2, giving d(s1', s2') + 1
           - We know d(s1', s2') >= |s2'| - |s1'| by IH
           - If |s2'| > |s1'|, then d(s1', c2::s2') must account for the extra character
           - At minimum, d(s1', c2::s2') >= |c2::s2'| - |s1'| - 0 = S|s2'| - |s1'| >= |s2'| - |s1'|

           Let's use a simpler fact: since any distance is non-negative, and we're adding 1,
           we just need to show that the base distances satisfy bounds. *)

        (* min3 a b c >= k iff a >= k /\ b >= k /\ c >= k *)
        (* We'll show each branch individually *)
        unfold min3.

        (* Branch 1: lev_distance s1' (c2 :: s2') + 1 >= length s2' - length s1' *)
        assert (H_br1: lev_distance s1' (c2 :: s2') + 1 >= length s2' - length s1').
        { apply Nat.leb_le in E_len.
          assert (H_case: length s1' = length s2' \/ length s1' < length s2') by lia.
          destruct H_case as [H_eq | H_lt].
          - (* |s1'| = |s2'|, so bound is 0 *)
            rewrite H_eq. simpl. lia.
          - (* |s1'| < |s2'|, so |s2'| - |s1'| >= 1 *)
            (* We know |c2::s2'| = S|s2'| and |s1'| < |s2'| *)
            (* So ||c2::s2'| - |s1'|| = S|s2'| - |s1'| *)
            assert (H_IH': lev_distance s1' (c2 :: s2') >= abs_diff (length s1') (S (length s2'))).
            { apply IHs1. }
            unfold abs_diff in H_IH'.
            assert (H_cmp: length s1' <=? S (length s2') = true).
            { apply Nat.leb_le. lia. }
            rewrite H_cmp in H_IH'.
            (* Now H_IH': d(s1', c2::s2') >= S|s2'| - |s1'| *)
            (* We need: d(s1', c2::s2') + 1 >= |s2'| - |s1'| *)
            (* Since |s1'| < |s2'|, we have S|s2'| - |s1'| = 1 + |s2'| - |s1'| *)
            apply Nat.leb_le in E_len.
            lia. }

        (* Branch 2: lev_distance (c1 :: s1') s2' + 1 >= length s2' - length s1' *)
        assert (H_br2: lev_distance (c1 :: s1') s2' + 1 >= length s2' - length s1').
        { (* Observe that d(c1::s1', s2') >= d(s1', s2') when we can delete c1 *)
          (* By definition: d(c1::s1', s2') = min3(d(s1', s2')+1, d(c1::s1', [])+1, d(s1', [])+subst) *)
          (* Actually, by definition: d(c1::s1', s2') = min3(...) which includes d(s1', s2')+subst as one branch *)
          (* So d(c1::s1', s2') <= d(s1', s2') + 1 *)
          (* But we need a lower bound. Note that one of the branches is d(s1', s2') + 0or1 *)
          (* The substitution branch gives d(s1', s2') + subst_cost c1 c_first_of_s2 *)
          (* Actually, let's use: to go from c1::s1' to s2', we can delete c1 (cost 1) then go s1' to s2' *)
          (* So d(c1::s1', s2') <= d(s1', s2') + 1 *)
          (* But we need >=, not <=! *)
          (*
          Hmm, the key insight: d(c1::s1', s2') by the recursive definition considers deleting c1,
          which gives branch d(s1', s2') + 1. Since lev_distance returns the MIN, we have:
            d(c1::s1', s2') <= d(s1', s2') + 1
          But for a LOWER bound, we need to think differently.

          Alternative: Since |s1'| <= |s2'|, adding c1 makes |c1::s1'| = S|s1'|.
          Case 1: S|s1'| <= |s2'|. Then|s2'| - |s1'| >= 1.
                  Since any edit distance >= 0, d(c1::s1', s2') + 1 >= 1.
                  If |s2'| - |s1'| = 1, we're done.
                  If |s2'| - |s1'| > 1, we need d(c1::s1', s2') + 1 >= |s2'| - |s1'| > 1,
                  so d(c1::s1', s2') >= |s2'| - |s1'| - 1 = |s2'| - S|s1'|.

          Actually, observe: transforming c1::s1' (length S|s1'|) to s2' (length |s2'|)
          requires at least ||s2'| - S|s1'|| edits (intuitive lower bound).
          When S|s1'| < |s2'|, this is |s2'| - S|s1'| = (|s2'| - |s1'|) - 1.
          So d(c1::s1', s2') >= |s2'| - |s1'| - 1, thus d + 1 >= |s2'| - |s1'|.

          But I haven't proven this "intuitive lower bound" - that's exactly the lemma I'm proving!
          This is circular.

          Solution: Use well-founded induction on length s1 + length s2.
          But changing induction strategy now is too disruptive.

          Pragmatic solution: Prove a helper lemma about deletion.
          OR: Observe that the one-char deletion bound is easy to prove directly.
          *)

          (* Direct approach: d(c1::s1', s2') can delete c1 to get d(s1', s2'), costing 1 *)
          (* So d(c1::s1', s2') is the min of several options including "delete c1" *)
          (* This means d(c1::s1', s2') <= d(s1', s2') + 1 *)
          (* But I need a lower bound! The issue is that the MIN could be much smaller. *)

          (* Let me try a different approach: use the contrapositive of upper bound *)
          (* Actually no, upper bound doesn't help with lower bound. *)

          (* Key realization: I can use the IH on s1' to get d(s1', s2') >= |s2'| - |s1'| *)
          (* Then observe that deleting c1 from c1::s1' costs 1, so: *)
          (* d(c1::s1', s2') + 1 >= d(via delete c1) + 1 = (d(s1', s2') + 1) + 1 = d(s1', s2') + 2 *)
          (* But this gives >= |s2'| - |s1'| + 2, which is too strong (>=, not what we want) *)

          (* Wait, deleting c1 is ONE way to transform, so d(c1::s1', s2') <= d(s1', s2') + 1 *)
          (* That's an upper bound on d(c1::s1', s2'), not useful for proving >= *)

          (* New approach: split by whether s2' is empty or not *)
          (* But wait - E_len refers to s2', and if I destruct it the hypothesis becomes invalid *)
          (* Better: just admit the whole branch 2, we'll fix with well-founded recursion *)
          (*
          The issue is circular: to prove d(c1::s1', s2') >= |s2'| - |s1'| when |s1'| < |s2'|,
          we'd need the very lemma we're proving (for strings of total length |c1::s1'| + |s2'|).
          Simple structural induction on s1 is insufficient.

          SOLUTION: Admit Branch 2 for now. Will reprove entire lemma using well-founded induction
          on (length s1 + length s2) later.
          *)
          admit.
        }

        (* Now combine all three branches *)
        (* Goal: min3 a b c >= k, where min3 a b c = min (min a b) c *)
        (* We've shown a >= k (H_br1), b >= k (H_br2), c >= k (H_br3) *)
        (* Therefore min (min a b) c >= k *)
        unfold min3.
        (* The min of values all >= k is also >= k *)
        (* min3 a b c = min a (min b c) *)
        assert (H: forall x y z k, x >= k -> y >= k -> z >= k -> Nat.min x (Nat.min y z) >= k).
        { intros x y z k Hx Hy Hz.
          apply Nat.min_case; [assumption | apply Nat.min_case; assumption]. }
        apply H; [exact H_br1 | exact H_br2 | exact H_br3].

      * (* |s1'| > |s2'|, so abs_diff = |s1'| - |s2'| *)
        (* This case is symmetric to the previous one *)
        (* By symmetry: d(c1::s1', c2::s2') = d(c2::s2', c1::s1') *)
        (* The proof structure is identical, just with roles reversed *)
        (* Since the previous case had Branch 2 admitted due to circularity, *)
        (* this case will have the same issue *)
        (* For now, admit the entire second case - will reprove with well-founded induction *)
        admit.
Admitted.
*)
*)

(* ========================================================================== *)
(* TRACE-BASED PROOF OF TRIANGLE INEQUALITY                                   *)
(* Based on Wagner & Fischer (1974) "The String-to-String Correction Problem" *)
(* ========================================================================== *)

(**
   Trace Abstraction:

   A trace from string A to B is a formalization of how an edit sequence transforms
   A into B, abstracting away the order of operations and focusing on the correspondence
   between character positions.

   Intuitively, a trace is a set of "matching lines" connecting position i in A to
   position j in B, where:
   - Each position is touched by at most one line
   - Lines don't cross (order-preserving)
   - Untouched positions represent insertions/deletions

   Reference: Wagner & Fischer (1974), Section 3 "Traces"
*)

(** A trace is represented as a list of pairs (i, j) where 1 <= i <= |A|, 1 <= j <= |B| *)
Definition Trace (A B : list Char) := list (nat * nat).

(** Check if a pair is valid for given string lengths *)
Definition valid_pair (lenA lenB : nat) (p : nat * nat) : bool :=
  let (i, j) := p in
  (1 <=? i) && (i <=? lenA) && (1 <=? j) && (j <=? lenB).

(** Check if two pairs are compatible (don't violate trace conditions) *)
Definition compatible_pairs (p1 p2 : nat * nat) : bool :=
  let '(i1, j1) := p1 in
  let '(i2, j2) := p2 in
  (* Different positions must not touch same indices, and must preserve order *)
  if (i1 =? i2) && (j1 =? j2) then true  (* same pair *)
  else if (i1 =? i2) || (j1 =? j2) then false  (* touch same position *)
  else
    (* Preserve order: i1 < i2 iff j1 < j2 (lines don't cross) *)
    if i1 <? i2 then j1 <? j2 else j2 <? j1.

(** Check if a list of pairs forms a valid trace *)
Fixpoint is_valid_trace_aux (pairs : list (nat * nat)) : bool :=
  match pairs with
  | [] => true
  | p :: ps =>
      (forallb (compatible_pairs p) ps) && is_valid_trace_aux ps
  end.

Definition is_valid_trace (A B : list Char) (T : Trace A B) : bool :=
  (forallb (valid_pair (length A) (length B)) T) && is_valid_trace_aux T.

(** Calculate which positions are touched by the trace *)
Fixpoint touched_in_A (A B : list Char) (T : Trace A B) : list nat :=
  match T with
  | [] => []
  | (i, _) :: rest => i :: touched_in_A A B rest
  end.

Fixpoint touched_in_B (A B : list Char) (T : Trace A B) : list nat :=
  match T with
  | [] => []
  | (_, j) :: rest => j :: touched_in_B A B rest
  end.

(** Cost of a trace according to Wagner-Fischer definition *)
Definition trace_cost (A B : list Char) (T : Trace A B) : nat :=
  (* Cost of change operations for matched pairs *)
  let change_cost := fold_left (fun acc p =>
    let '(i, j) := p in
    acc + subst_cost (nth (i-1) A default_char) (nth (j-1) B default_char)
  ) T 0 in

  (* Cost of deletions (positions in A not touched) *)
  let delete_cost := length A - length (touched_in_A A B T) in

  (* Cost of insertions (positions in B not touched) *)
  let insert_cost := length B - length (touched_in_B A B T) in

  change_cost + delete_cost + insert_cost.

(**
   Trace Composition (Wagner-Fischer, page 3):

   If T1 is a trace from A to B and T2 is a trace from B to C,
   then T1 ∘ T2 is defined as the trace from A to C where:

   (i, k) ∈ T1 ∘ T2  iff  ∃j such that (i,j) ∈ T1 and (j,k) ∈ T2

   This represents composing the transformations: A → B → C becomes A → C
*)
Definition compose_trace {A B C : list Char} (T1 : Trace A B) (T2 : Trace B C) : Trace A C :=
  fold_left (fun acc p1 =>
    let '(i, j) := p1 in
    (* Find all pairs (j, k) in T2 where first component matches j *)
    let matches := filter (fun p2 => let '(j2, k) := p2 in j =? j2) T2 in
    (* Add (i, k) for each match *)
    fold_left (fun acc2 p2 =>
      let '(_, k) := p2 in
      (i, k) :: acc2
    ) matches acc
  ) T1 [].

(** Helper lemmas for compose_trace_preserves_validity *)

(**
   Helper: Membership in fold_left for the inner fold pattern used in compose_trace.

   When we fold over matches to build pairs (i,k), an element appears in the result
   if it was already in the accumulator or it's one of the newly added pairs.
*)
Lemma In_fold_left_cons_pairs :
  forall (i : nat) (matches : list (nat * nat)) (acc : list (nat * nat)) (k : nat),
    In (i, k) (fold_left (fun acc2 p2 => let '(_, k') := p2 in (i, k') :: acc2) matches acc) <->
    In (i, k) acc \/ exists j, In (j, k) matches.
Proof.
  intros i matches.
  induction matches as [| [j' k'] matches' IH]; intros acc k.
  - (* Base case: matches = [] *)
    simpl.
    split; intro H.
    + left. exact H.
    + destruct H as [H | [j H]].
      * exact H.
      * contradiction.
  - (* Inductive case: matches = (j', k') :: matches' *)
    simpl.
    rewrite IH.
    split; intro H.
    + destruct H as [H | [j H]].
      * (* (i,k) was in the new acc after adding (i,k') *)
        simpl in H.
        destruct H as [H | H].
        -- (* (i,k) = (i,k') *)
           inversion H; subst.
           right. exists j'. left. reflexivity.
        -- (* (i,k) was in original acc *)
           left. exact H.
      * (* exists j witness in matches' *)
        right. exists j. right. exact H.
    + destruct H as [H | [j H]].
      * (* (i,k) in original acc *)
        left. simpl. right. exact H.
      * (* exists j witness in full matches *)
        simpl in H.
        destruct H as [H | H].
        -- (* j = j', k was paired with j' *)
           inversion H; subst.
           left. simpl. left. reflexivity.
        -- (* j witness is in matches' *)
           right. exists j. exact H.
Qed.

(**
   Helper: Connection between filter and membership.

   A pair (j,k) is in the filtered list iff it's in T2 and j matches the filter criterion.
*)
Lemma In_filter_eq :
  forall (j_target : nat) (T2 : list (nat * nat)) (j k : nat),
    In (j, k) (filter (fun p2 => let '(j2, _) := p2 in j_target =? j2) T2) <->
    In (j, k) T2 /\ j_target = j.
Proof.
  intros j_target T2 j k.
  rewrite filter_In.
  split; intro H.
  - destruct H as [H_in H_eq].
    simpl in H_eq.
    apply Nat.eqb_eq in H_eq.
    split; assumption.
  - destruct H as [H_in H_eq].
    split.
    + exact H_in.
    + simpl. apply Nat.eqb_eq. exact H_eq.
Qed.

(**
   Helper: The inner fold preserves membership from accumulator.

   Any pair in the accumulator remains in the result.
*)
Lemma In_fold_preserves_acc :
  forall (i' : nat) (matches acc : list (nat * nat)) (p : nat * nat),
    In p acc ->
    In p (fold_left (fun acc2 p2 => let '(_, k') := p2 in (i', k') :: acc2) matches acc).
Proof.
  intros i' matches.
  induction matches as [| [j_m k_m] matches' IH]; intros acc p H_in.
  - (* Base: matches = [] *)
    simpl. exact H_in.
  - (* Inductive: matches = (j_m, k_m) :: matches' *)
    simpl.
    apply IH.
    simpl. right. exact H_in.
Qed.

(**
   Helper: If i ≠ i', then pairs (i, k) in the fold result must have been in acc.

   The fold only adds pairs of form (i', k'), so pairs with a different first component
   must have come from the accumulator.
*)
Lemma In_fold_diff_first :
  forall (i i' : nat) (matches acc : list (nat * nat)) (k : nat),
    i <> i' ->
    In (i, k) (fold_left (fun acc2 p2 => let '(_, k') := p2 in (i', k') :: acc2) matches acc) ->
    In (i, k) acc.
Proof.
  intros i i' matches.
  induction matches as [| [j_m k_m] matches' IH]; intros acc k H_neq H_in.
  - (* Base: matches = [] *)
    simpl in H_in. exact H_in.
  - (* Inductive: matches = (j_m, k_m) :: matches' *)
    simpl in H_in.
    apply IH in H_in; [| exact H_neq].
    simpl in H_in.
    destruct H_in as [H_eq | H_in].
    + (* (i, k) = (i', k_m) - contradiction since i ≠ i' *)
      inversion H_eq; subst.
      exfalso. apply H_neq. reflexivity.
    + (* (i, k) was in original acc *)
      exact H_in.
Qed.

(**
   Helper: Membership in the outer fold_left of compose_trace.

   This lemma characterizes when a pair appears in the accumulating result
   of the composition fold operation.
*)
Lemma In_compose_trace_fold :
  forall (T1 : list (nat * nat)) (T2 : list (nat * nat)) (acc : list (nat * nat)) (i k : nat),
    In (i, k) (fold_left (fun acc' p1 =>
      let '(i', j) := p1 in
      let matches := filter (fun p2 => let '(j2, _) := p2 in j =? j2) T2 in
      fold_left (fun acc2 p2 => let '(_, k') := p2 in (i', k') :: acc2) matches acc'
    ) T1 acc) <->
    In (i, k) acc \/ exists j, In (i, j) T1 /\ In (j, k) T2.
Proof.
  intros T1 T2.
  induction T1 as [| [i' j'] T1' IH]; intros acc i k.
  - (* Base case: T1 = [] *)
    simpl.
    split; intro H.
    + left. exact H.
    + destruct H as [H | [j [H _]]].
      * exact H.
      * contradiction.
  - (* Inductive case: T1 = (i',j') :: T1' *)
    simpl.
    split; intro H.
    + (* Forward: membership in result -> witness or in acc *)
      rewrite IH in H.
      destruct H as [H | [j [H_in1 H_in2]]].
      * (* (i,k) is in the new accumulator after processing (i',j') *)
        (* Key insight: the inner fold ONLY adds pairs of form (i', k').
           So if In (i,k) holds in the result, either:
           - (i,k) was already in acc, OR
           - i = i' and k came from a match *)
        destruct (Nat.eq_dec i i') as [H_eq | H_neq].
        -- (* Case: i = i' *)
           subst i'.
           set (matches := filter (fun p2 : nat * nat => let '(j2, _) := p2 in j' =? j2) T2) in H.
           pose proof (In_fold_left_cons_pairs i matches acc k) as H_inner.
           rewrite H_inner in H. clear H_inner.
           destruct H as [H_acc | [j_m H_match]].
           ++ (* Was in acc *)
              left. exact H_acc.
           ++ (* Came from match *)
              unfold matches in H_match.
              rewrite In_filter_eq in H_match.
              destruct H_match as [H_in_T2 H_j_eq].
              subst j_m.
              (* We have (j', k) ∈ T2, and the pair (i, j') is in the current position of T1 *)
              right. exists j'. split.
              ** left. reflexivity.
              ** exact H_in_T2.
        -- (* Case: i ≠ i' *)
           (* The fold only adds pairs (i', k'), so In (i, k) must have been in acc *)
           set (matches := filter (fun p2 : nat * nat => let '(j2, _) := p2 in j' =? j2) T2) in H.
           apply In_fold_diff_first in H; [| exact H_neq].
           left. exact H.
      * (* There's a witness in T1' *)
        right. exists j. split.
        -- right. exact H_in1.
        -- exact H_in2.
    + (* Backward: witness or in acc -> membership in result *)
      rewrite IH.
      destruct H as [H | [j [H_in1 H_in2]]].
      * (* Was in original acc *)
        (* Since (i,k) is in acc, it remains in the fold result *)
        set (matches := filter (fun p2 : nat * nat => let '(j2, _) := p2 in j' =? j2) T2).
        left.
        apply In_fold_preserves_acc.
        exact H.
      * (* There's a witness *)
        simpl in H_in1.
        destruct H_in1 as [H_eq | H_in1].
        -- (* Witness is (i',j') itself *)
           inversion H_eq; subst.
           (* Now i=i', j=j', and we have (j',k) ∈ T2 *)
           (* We need to show (i,k) is in fold result after processing (i,j') *)
           (* The filter will find (j',k) in T2, and fold will add (i,k) *)
           set (matches := filter (fun p2 : nat * nat => let '(j2, _) := p2 in j =? j2) T2).
           pose proof (In_fold_left_cons_pairs i matches acc k) as H_inner.
           left.
           rewrite H_inner.
           right. exists j.
           unfold matches.
           rewrite In_filter_eq.
           split; [exact H_in2 | reflexivity].
        -- (* Witness is in T1' *)
           right. exists j. split; assumption.
Qed.

(**
   Characterization of membership in composed trace.

   A pair (i,k) appears in the composed trace iff there exists some j
   such that (i,j) is in T1 and (j,k) is in T2.
*)
Lemma In_compose_trace :
  forall (A B C : list Char) (T1 : Trace A B) (T2 : Trace B C) (i k : nat),
    In (i, k) (compose_trace T1 T2) <->
    exists j, In (i, j) T1 /\ In (j, k) T2.
Proof.
  intros A B C T1 T2 i k.
  unfold compose_trace.
  rewrite In_compose_trace_fold with (acc := []).
  split; intro H.
  - (* Forward direction *)
    destruct H as [H | H].
    + (* In empty list - contradiction *)
      contradiction.
    + (* Exists witness *)
      exact H.
  - (* Backward direction *)
    right. exact H.
Qed.

(** Helper lemmas for compose_trace_preserves_validity *)

(**
   Valid pairs compose transitively.

   If (i,j) is valid for strings of length |A| and |B|,
   and (j,k) is valid for strings of length |B| and |C|,
   then (i,k) is valid for strings of length |A| and |C|.
*)
Lemma valid_pair_compose :
  forall (lenA lenB lenC : nat) (i j k : nat),
    valid_pair lenA lenB (i, j) = true ->
    valid_pair lenB lenC (j, k) = true ->
    valid_pair lenA lenC (i, k) = true.
Proof.
  intros lenA lenB lenC i j k H1 H2.
  unfold valid_pair in *.
  simpl in *.
  (* Structure after unfolding:
     H1: (1 <=? i) && (i <=? lenA) && (1 <=? j) && (j <=? lenB) = true
     H2: (1 <=? j) && (j <=? lenB) && (1 <=? k) && (k <=? lenC) = true
     Goal: (1 <=? i) && (i <=? lenA) && (1 <=? k) && (k <=? lenC) = true
  *)

  (* Extract bounds from H1: need (1 <=? i) and (i <=? lenA) *)
  apply andb_true_iff in H1 as [H1_left H1_jB].
  apply andb_true_iff in H1_left as [H1_left2 H1_jlow].
  apply andb_true_iff in H1_left2 as [H1_ilow H1_ihigh].

  (* Extract bounds from H2: need (1 <=? k) and (k <=? lenC) *)
  apply andb_true_iff in H2 as [H2_left H2_kC].
  apply andb_true_iff in H2_left as [H2_left2 H2_klow].
  apply andb_true_iff in H2_left2 as [H2_jlow H2_jB].

  (* Construct the result: (1 <=? i) && (i <=? lenA) && (1 <=? k) && (k <=? lenC) *)
  apply andb_true_intro. split.
  - apply andb_true_intro. split.
    + apply andb_true_intro. split.
      * exact H1_ilow.
      * exact H1_ihigh.
    + exact H2_klow.
  - exact H2_kC.
Qed.

(** * Infrastructure for Trace Validity Preservation *)

(**
   Extract order preservation from compatible_pairs.

   If two pairs are compatible and have different components, then their
   first and second components preserve the same order.
*)
Lemma compatible_pairs_order :
  forall (i1 j1 i2 j2 : nat),
    i1 <> i2 ->
    j1 <> j2 ->
    compatible_pairs (i1, j1) (i2, j2) = true ->
    (i1 < i2 <-> j1 < j2).
Proof.
  intros i1 j1 i2 j2 H_i_neq H_j_neq H_compat.
  unfold compatible_pairs in H_compat.
  simpl in H_compat.

  (* The compatible_pairs definition checks:
     if i1 =? i2 && j1 =? j2 then true  (rejected by H_i_neq, H_j_neq)
     else if i1 =? i2 || j1 =? j2 then false  (must be false for H_compat to be true)
     else if i1 <? i2 then j1 <? j2 else j2 <? j1
  *)

  (* Case analysis based on the structure of compatible_pairs *)
  destruct (i1 =? i2) eqn:H_i_eq.
  - (* i1 = i2 - contradiction *)
    apply Nat.eqb_eq in H_i_eq.
    exfalso. apply H_i_neq. exact H_i_eq.
  - (* i1 <> i2 *)
    destruct (j1 =? j2) eqn:H_j_eq.
    + (* j1 = j2 - contradiction *)
      apply Nat.eqb_eq in H_j_eq.
      exfalso. apply H_j_neq. exact H_j_eq.
    + (* j1 <> j2 *)
      (* Now we're in the third case: if i1 <? i2 then j1 <? j2 else j2 <? j1 *)
      simpl in H_compat.
      destruct (i1 <? i2) eqn:H_i_ltb.
      * (* i1 < i2 *)
        apply Nat.ltb_lt in H_i_ltb.
        apply Nat.ltb_lt in H_compat.
        split; intro; assumption.
      * (* i1 >= i2, so i2 < i1 (since i1 <> i2) *)
        apply Nat.ltb_ge in H_i_ltb.
        apply Nat.ltb_lt in H_compat.
        assert (H_i2_lt: i2 < i1).
        { apply Nat.eqb_neq in H_i_eq. lia. }
        split; intro H; exfalso; lia.
Qed.

(**
   Valid traces have unique first components.

   If a valid trace contains two pairs with the same first component,
   they must have the same second component (i.e., each position in the
   source can match at most one position in the target).
*)
Lemma valid_trace_unique_first :
  forall (T : list (nat * nat)) (i j1 j2 : nat),
    is_valid_trace_aux T = true ->
    In (i, j1) T ->
    In (i, j2) T ->
    j1 = j2.
Proof.
  intros T i j1 j2 H_valid H_in1 H_in2.
  induction T as [| [i' j'] T' IH].
  - (* Base case: T = [] *)
    contradiction.
  - (* Inductive case: T = (i', j') :: T' *)
    simpl in H_valid.
    apply andb_true_iff in H_valid as [H_forall H_valid'].

    simpl in H_in1, H_in2.
    destruct H_in1 as [H_eq1 | H_in1]; destruct H_in2 as [H_eq2 | H_in2].

    + (* (i, j1) = (i', j') and (i, j2) = (i', j') *)
      inversion H_eq1; inversion H_eq2; subst.
      reflexivity.

    + (* (i, j1) = (i', j') and (i, j2) ∈ T' *)
      inversion H_eq1; subst.
      clear H_eq1.
      (* Use compatibility: (i, j1) must be compatible with all pairs in T' *)
      rewrite forallb_forall in H_forall.
      specialize (H_forall (i, j2) H_in2).
      unfold compatible_pairs in H_forall.
      simpl in H_forall.
      (* Check if i =? i and j1 =? j2 *)
      rewrite Nat.eqb_refl in H_forall.
      simpl in H_forall.
      destruct (j1 =? j2) eqn:H_j_eq.
      * (* j1 = j2 *)
        apply Nat.eqb_eq in H_j_eq.
        exact H_j_eq.
      * (* j1 <> j2, but (i =? i) || (j1 =? j2) = true, making compatible_pairs false *)
        (* The definition says: if i1=i2 || j1=j2 then false (when not both equal) *)
        (* We have i=i (true) and j1≠j2, so the orb is true, result should be false *)
        discriminate H_forall.

    + (* (i, j1) ∈ T' and (i, j2) = (i', j') *)
      inversion H_eq2; subst.
      clear H_eq2.
      (* Similar to previous case, symmetric *)
      rewrite forallb_forall in H_forall.
      specialize (H_forall (i, j1) H_in1).
      unfold compatible_pairs in H_forall.
      simpl in H_forall.
      rewrite Nat.eqb_refl in H_forall.
      simpl in H_forall.
      destruct (j2 =? j1) eqn:H_j_eq.
      * apply Nat.eqb_eq in H_j_eq.
        symmetry. exact H_j_eq.
      * discriminate H_forall.

    + (* Both (i, j1) ∈ T' and (i, j2) ∈ T' *)
      apply IH; assumption.
Qed.

(**
   Valid traces have unique second components (symmetric version).

   If a valid trace contains two pairs with the same second component,
   they must have the same first component (i.e., each position in the
   target can be matched by at most one position in the source).
*)
Lemma valid_trace_unique_second :
  forall (T : list (nat * nat)) (i1 i2 j : nat),
    is_valid_trace_aux T = true ->
    In (i1, j) T ->
    In (i2, j) T ->
    i1 = i2.
Proof.
  intros T i1 i2 j H_valid H_in1 H_in2.
  induction T as [| [i' j'] T' IH].
  - (* Base case: T = [] *)
    contradiction.
  - (* Inductive case: T = (i', j') :: T' *)
    simpl in H_valid.
    apply andb_true_iff in H_valid as [H_forall H_valid'].

    simpl in H_in1, H_in2.
    destruct H_in1 as [H_eq1 | H_in1]; destruct H_in2 as [H_eq2 | H_in2].

    + (* (i1, j) = (i', j') and (i2, j) = (i', j') *)
      inversion H_eq1; inversion H_eq2; subst.
      reflexivity.

    + (* (i1, j) = (i', j') and (i2, j) ∈ T' *)
      inversion H_eq1; subst.
      clear H_eq1.
      (* Use compatibility: (i1, j) must be compatible with all pairs in T' *)
      rewrite forallb_forall in H_forall.
      specialize (H_forall (i2, j) H_in2).
      unfold compatible_pairs in H_forall.
      simpl in H_forall.
      (* Check if i1 =? i2 and j =? j *)
      destruct (i1 =? i2) eqn:H_i_eq.
      * (* i1 = i2 *)
        apply Nat.eqb_eq in H_i_eq.
        exact H_i_eq.
      * (* i1 <> i2, but j = j, so the orb (i1 =? i2) || (j =? j) = true *)
        rewrite Nat.eqb_refl in H_forall.
        simpl in H_forall.
        discriminate H_forall.

    + (* (i1, j) ∈ T' and (i2, j) = (i', j') *)
      inversion H_eq2; subst.
      clear H_eq2.
      (* Symmetric *)
      rewrite forallb_forall in H_forall.
      specialize (H_forall (i1, j) H_in1).
      unfold compatible_pairs in H_forall.
      simpl in H_forall.
      destruct (i2 =? i1) eqn:H_i_eq.
      * apply Nat.eqb_eq in H_i_eq.
        symmetry. exact H_i_eq.
      * rewrite Nat.eqb_refl in H_forall.
        simpl in H_forall.
        discriminate H_forall.

    + (* Both (i1, j) ∈ T' and (i2, j) ∈ T' *)
      apply IH; assumption.
Qed.

(**
   Order preservation in valid traces.

   If two distinct pairs are in a valid trace, their first and second
   components preserve the same ordering relationship.
*)
Lemma valid_trace_order_preserved :
  forall (T : list (nat * nat)) (i1 j1 i2 j2 : nat),
    is_valid_trace_aux T = true ->
    In (i1, j1) T ->
    In (i2, j2) T ->
    i1 <> i2 ->
    (i1 < i2 <-> j1 < j2).
Proof.
  intros T i1 j1 i2 j2 H_valid H_in1 H_in2 H_neq.

  (* First, prove that j1 <> j2 *)
  assert (H_j_neq: j1 <> j2).
  {
    intro H_j_eq.
    subst j2.
    (* If j1 = j2, then by uniqueness of second components, i1 = i2 *)
    assert (H_eq: i1 = i2).
    { apply (valid_trace_unique_second T i1 i2 j1 H_valid H_in1 H_in2). }
    contradiction.
  }

  (* Now extract compatibility from the valid trace *)
  induction T as [| [i' j'] T' IH].
  - (* Base: T = [] *)
    contradiction.
  - (* Inductive: T = (i', j') :: T' *)
    simpl in H_valid.
    apply andb_true_iff in H_valid as [H_forall H_valid'].

    simpl in H_in1, H_in2.
    destruct H_in1 as [H_eq1 | H_in1]; destruct H_in2 as [H_eq2 | H_in2].

    + (* Both equal (i', j') - contradiction with i1 <> i2 *)
      inversion H_eq1; inversion H_eq2; subst.
      exfalso. apply H_neq. reflexivity.

    + (* (i1, j1) = (i', j') and (i2, j2) ∈ T' *)
      inversion H_eq1; subst.
      clear H_eq1.
      (* Apply compatibility *)
      rewrite forallb_forall in H_forall.
      specialize (H_forall (i2, j2) H_in2).
      apply compatible_pairs_order; assumption.

    + (* (i1, j1) ∈ T' and (i2, j2) = (i', j') *)
      inversion H_eq2; subst.
      clear H_eq2.
      (* Apply compatibility - compatible_pairs (i2, j2) (i1, j1) *)
      rewrite forallb_forall in H_forall.
      specialize (H_forall (i1, j1) H_in1).
      (* Use compatible_pairs_order with swapped arguments *)
      assert (H_neq_sym: i2 <> i1).
      { intro H_eq. symmetry in H_eq. contradiction. }
      assert (H_j_neq_sym: j2 <> j1).
      { intro H_eq. symmetry in H_eq. contradiction. }
      apply compatible_pairs_order in H_forall; [| exact H_neq_sym | exact H_j_neq_sym].
      (* H_forall now gives us: i2 < i1 <-> j2 < j1 *)
      (* We need: i1 < i2 <-> j1 < j2, which is the contrapositive *)
      split; intro H.
      * (* i1 < i2 -> j1 < j2 *)
        assert (H_not_i2_lt: ~ (i2 < i1)).
        { lia. }
        assert (H_not_j2_lt: ~ (j2 < j1)).
        { intro H_j2_lt. apply H_not_i2_lt. apply H_forall. exact H_j2_lt. }
        lia.
      * (* j1 < j2 -> i1 < i2 *)
        assert (H_not_j2_lt: ~ (j2 < j1)).
        { lia. }
        assert (H_not_i2_lt: ~ (i2 < i1)).
        { intro H_i2_lt. apply H_not_j2_lt. apply H_forall. exact H_i2_lt. }
        lia.

    + (* Both in T' *)
      apply IH; assumption.
Qed.

(** * Helper Lemmas for Trace Validity Preservation *)

(**
   Extract pairwise compatibility from valid trace.

   If a trace is valid (is_valid_trace_aux = true), then any two pairs
   in the trace are compatible with each other.
*)
Lemma is_valid_trace_aux_In_compatible :
  forall (T : list (nat * nat)) (p1 p2 : nat * nat),
    is_valid_trace_aux T = true ->
    In p1 T ->
    In p2 T ->
    compatible_pairs p1 p2 = true.
Proof.
  intros T p1 p2 H_valid H_in1 H_in2.
  induction T as [| p T' IH].
  - (* Base: T = [] *)
    contradiction.
  - (* Inductive: T = p :: T' *)
    simpl in H_valid.
    apply andb_true_iff in H_valid as [H_forall H_valid'].

    simpl in H_in1, H_in2.
    destruct H_in1 as [H_eq1 | H_in1]; destruct H_in2 as [H_eq2 | H_in2].

    + (* p1 = p and p2 = p *)
      subst p1 p2.
      unfold compatible_pairs.
      destruct p as [i j].
      simpl.
      rewrite Nat.eqb_refl.
      rewrite Nat.eqb_refl.
      reflexivity.

    + (* p1 = p and p2 ∈ T' *)
      subst p1.
      rewrite forallb_forall in H_forall.
      apply H_forall.
      exact H_in2.

    + (* p1 ∈ T' and p2 = p *)
      subst p2.
      rewrite forallb_forall in H_forall.
      (* Need to use symmetry of compatible_pairs *)
      assert (H_compat: compatible_pairs p p1 = true).
      { apply H_forall. exact H_in1. }
      (* compatible_pairs is symmetric *)
      unfold compatible_pairs in *.
      destruct p as [i_p j_p].
      destruct p1 as [i1 j1].
      simpl in *.
      destruct (i_p =? i1) eqn:H_i_eq; destruct (j_p =? j1) eqn:H_j_eq.
      * (* Both equal - use symmetry of =? *)
        apply Nat.eqb_eq in H_i_eq, H_j_eq.
        subst i1 j1.
        rewrite Nat.eqb_refl.
        rewrite Nat.eqb_refl.
        reflexivity.
      * simpl in H_compat. discriminate.
      * simpl in H_compat. discriminate.
      * simpl in H_compat.
        (* Need to show compatible_pairs (i1,j1) (i_p,j_p) given compatible_pairs (i_p,j_p) (i1,j1) *)
        (* Both i and j are different, so check order *)
        destruct (i1 =? i_p) eqn:H_i_eq2.
        -- (* i1 = i_p contradicts i_p <> i1 *)
           apply Nat.eqb_eq in H_i_eq2.
           apply Nat.eqb_neq in H_i_eq.
           exfalso. apply H_i_eq. symmetry. exact H_i_eq2.
        -- destruct (j1 =? j_p) eqn:H_j_eq2.
           ++ (* j1 = j_p contradicts j_p <> j1 *)
              apply Nat.eqb_eq in H_j_eq2.
              apply Nat.eqb_neq in H_j_eq.
              exfalso. apply H_j_eq. symmetry. exact H_j_eq2.
           ++ (* Both different - use order reversal *)
              simpl.
              destruct (i_p <? i1) eqn:H_i_lt.
              ** (* i_p < i1, so we need i1 > i_p, which means i_p < i1, and j1 > j_p *)
                 apply Nat.ltb_lt in H_i_lt.
                 apply Nat.ltb_lt in H_compat.
                 (* Goal: (if i1 <? i_p then j1 <? j_p else j_p <? j1) = true *)
                 (* Since i_p < i1, we have ~(i1 < i_p), so the else branch applies *)
                 destruct (i1 <? i_p) eqn:H_i1_lt.
                 --- apply Nat.ltb_lt in H_i1_lt. exfalso. lia.
                 --- (* else branch: j_p <? j1 *)
                     apply Nat.ltb_lt. exact H_compat.
              ** (* i_p >= i1 and i_p <> i1, so i1 < i_p, and j1 < j_p *)
                 apply Nat.ltb_ge in H_i_lt.
                 apply Nat.ltb_lt in H_compat.
                 (* Since i1 < i_p, the then branch applies: need j1 < j_p *)
                 assert (H_i1_lt: i1 < i_p).
                 { apply Nat.eqb_neq in H_i_eq. lia. }
                 apply Nat.ltb_lt in H_i1_lt.
                 rewrite H_i1_lt.
                 apply Nat.ltb_lt. exact H_compat.

    + (* p1 ∈ T' and p2 ∈ T' *)
      apply IH; assumption.
Qed.

(**
   Build valid trace from pairwise compatibility.

   If all pairs in a list are pairwise compatible, then the list
   satisfies is_valid_trace_aux.
*)
Lemma is_valid_trace_aux_from_pairwise :
  forall (T : list (nat * nat)),
    (forall p1 p2, In p1 T -> In p2 T -> compatible_pairs p1 p2 = true) ->
    is_valid_trace_aux T = true.
Proof.
  induction T as [| p ps IH].
  - (* Base: T = [] *)
    intro H_pairwise.
    reflexivity.
  - (* Inductive: T = p :: ps *)
    intro H_pairwise.
    simpl.
    apply andb_true_iff.
    split.
    + (* forallb (compatible_pairs p) ps = true *)
      apply forallb_forall.
      intros p' H_in_ps.
      apply H_pairwise.
      * left. reflexivity.
      * right. exact H_in_ps.
    + (* is_valid_trace_aux ps = true *)
      apply IH.
      intros p1 p2 H_in1 H_in2.
      apply H_pairwise.
      * right. exact H_in1.
      * right. exact H_in2.
Qed.

(**
   Compatible pairs compose transitively.

   If two pairs from a composed trace have witnesses in the original traces,
   then they are compatible (order-preserving, no crossing).

   Key insight: If (i₁,j₁) and (i₂,j₂) are compatible in T1,
   and (j₁,k₁) and (j₂,k₂) are compatible in T2,
   then (i₁,k₁) and (i₂,k₂) are compatible (transitivity of order).
*)
Lemma compatible_pairs_compose :
  forall (T1 T2 : list (nat * nat)) (i1 j1 k1 i2 j2 k2 : nat),
    is_valid_trace_aux T1 = true ->
    is_valid_trace_aux T2 = true ->
    In (i1, j1) T1 ->
    In (i2, j2) T1 ->
    In (j1, k1) T2 ->
    In (j2, k2) T2 ->
    compatible_pairs (i1, k1) (i2, k2) = true.
Proof.
  intros T1 T2 i1 j1 k1 i2 j2 k2 H_valid1 H_valid2 H_in11 H_in12 H_in21 H_in22.
  unfold compatible_pairs.
  simpl.
  (* Case analysis on whether the pairs are the same *)
  destruct (Nat.eq_dec i1 i2) as [H_i_eq | H_i_neq].
  - (* i1 = i2 *)
    subst i2.
    destruct (Nat.eq_dec k1 k2) as [H_k_eq | H_k_neq].
    + (* k1 = k2: pairs are equal *)
      subst k2.
      rewrite Nat.eqb_refl.
      rewrite Nat.eqb_refl.
      reflexivity.
    + (* k1 ≠ k2 but i1 = i2 *)
      (* Since T1 is valid and contains (i1,j1) and (i1,j2), we must have j1 = j2 *)
      assert (H_j_eq: j1 = j2).
      { apply (valid_trace_unique_first T1 i1 j1 j2 H_valid1 H_in11 H_in12). }
      subst j2.
      (* Now T2 contains (j1,k1) and (j1,k2) with k1 ≠ k2 *)
      (* By uniqueness of first components in T2, this is impossible *)
      assert (H_k_eq: k1 = k2).
      { apply (valid_trace_unique_first T2 j1 k1 k2 H_valid2 H_in21 H_in22). }
      (* But we have k1 ≠ k2, contradiction *)
      exfalso. apply H_k_neq. exact H_k_eq.
  - (* i1 ≠ i2 *)
    destruct (Nat.eq_dec k1 k2) as [H_k_eq | H_k_neq].
    + (* k1 = k2 but i1 ≠ i2 *)
      (* Since T2 is valid and contains (j1,k1) and (j2,k2) with k1=k2, we must have j1 = j2 *)
      subst k2.
      assert (H_j_eq: j1 = j2).
      { apply (valid_trace_unique_second T2 j1 j2 k1 H_valid2 H_in21 H_in22). }
      subst j2.
      (* Now T1 contains (i1,j1) and (i2,j1) with i1 ≠ i2 *)
      (* By uniqueness of second components in T1, this is impossible *)
      assert (H_i_eq: i1 = i2).
      { apply (valid_trace_unique_second T1 i1 i2 j1 H_valid1 H_in11 H_in12). }
      (* But we have i1 ≠ i2, contradiction *)
      exfalso. apply H_i_neq. exact H_i_eq.
    + (* i1 ≠ i2 and k1 ≠ k2 *)
      (* Show order preservation: i1 < i2 ⟺ k1 < k2 *)
      (* By transitivity through the intermediate string B *)

      (* Get order preservation for T1: i1 < i2 ⟺ j1 < j2 *)
      assert (H_order1: i1 < i2 <-> j1 < j2).
      { apply (valid_trace_order_preserved T1 i1 j1 i2 j2 H_valid1 H_in11 H_in12 H_i_neq). }

      (* Get order preservation for T2: j1 < j2 ⟺ k1 < k2 *)
      (* First check if j1 = j2 *)
      destruct (Nat.eq_dec j1 j2) as [H_j_eq | H_j_neq].
      * (* j1 = j2 - then from T1, we'd have i1 = i2, contradiction *)
        subst j2.
        assert (H_i_eq: i1 = i2).
        { apply (valid_trace_unique_second T1 i1 i2 j1 H_valid1 H_in11 H_in12). }
        exfalso. apply H_i_neq. exact H_i_eq.
      * (* j1 ≠ j2 *)
        assert (H_order2: j1 < j2 <-> k1 < k2).
        { apply (valid_trace_order_preserved T2 j1 k1 j2 k2 H_valid2 H_in21 H_in22 H_j_neq). }

        (* Combine the two: i1 < i2 ⟺ j1 < j2 ⟺ k1 < k2 *)
        (* This gives us i1 < i2 ⟺ k1 < k2 *)
        (* Work directly with the boolean conditions *)
        destruct (i1 =? i2) eqn:H_i_eqb.
        -- (* i1 = i2 - contradiction *)
           apply Nat.eqb_eq in H_i_eqb.
           exfalso. apply H_i_neq. exact H_i_eqb.
        -- (* i1 <> i2 *)
           destruct (k1 =? k2) eqn:H_k_eqb.
           ++ (* k1 = k2 - contradiction *)
              apply Nat.eqb_eq in H_k_eqb.
              exfalso. apply H_k_neq. exact H_k_eqb.
           ++ (* Both different, check order *)
              simpl.
              destruct (i1 <? i2) eqn:H_i_ltb.
              ** (* i1 < i2 *)
                 destruct (k1 <? k2) eqn:H_k_ltb.
                 --- (* k1 < k2 - both orders match, result true *)
                     reflexivity.
                 --- (* k1 >= k2 - orders don't match, contradiction *)
                     apply Nat.ltb_lt in H_i_ltb.
                     apply Nat.ltb_ge in H_k_ltb.
                     apply H_order1 in H_i_ltb as H_j_lt.
                     apply H_order2 in H_j_lt as H_k_lt.
                     exfalso. lia.
              ** (* i1 >= i2, so i2 < i1 (since i1 <> i2) *)
                 destruct (k1 <? k2) eqn:H_k_ltb.
                 --- (* k1 < k2 - orders don't match, contradiction *)
                     apply Nat.ltb_ge in H_i_ltb.
                     apply Nat.ltb_lt in H_k_ltb.
                     assert (H_j_lt: j1 < j2).
                     { apply H_order2. exact H_k_ltb. }
                     assert (H_i_lt: i1 < i2).
                     { apply H_order1. exact H_j_lt. }
                     exfalso. lia.
                 --- (* k1 >= k2, so k2 < k1 (since k1 <> k2) - both reversed, result is k2 <? k1 *)
                     (* The goal is (if i2 <? i1 then k2 <? k1 else k1 <? k2) = true *)
                     (* Since i1 >= i2 and i1 <> i2, we have i2 < i1 *)
                     apply Nat.ltb_ge in H_i_ltb.
                     apply Nat.ltb_ge in H_k_ltb.
                     assert (H_i2_lt: i2 < i1).
                     { apply Nat.eqb_neq in H_i_eqb. lia. }
                     (* We have i2 < i1, so we need to show k2 < k1 *)
                     (* From i2 < i1, we get j2 < j1 (contrapositive of H_order1) *)
                     assert (H_j2_lt: j2 < j1).
                     { destruct H_order1 as [H_fwd H_bwd].
                       assert (H_not_i_lt: ~ (i1 < i2)).
                       { lia. }
                       assert (H_not_j_lt: ~ (j1 < j2)).
                       { intro H_j_lt. apply H_not_i_lt. apply H_bwd. exact H_j_lt. }
                       lia. }
                     (* From j2 < j1, we get k2 < k1 (by H_order2 contrapositive) *)
                     assert (H_k2_lt: k2 < k1).
                     { destruct H_order2 as [H_fwd H_bwd].
                       assert (H_not_j_lt: ~ (j1 < j2)).
                       { lia. }
                       assert (H_not_k_lt: ~ (k1 < k2)).
                       { intro H_k_lt. apply H_not_j_lt. apply H_bwd. exact H_k_lt. }
                       lia. }
                     (* Now apply Nat.ltb_lt to convert k2 < k1 to k2 <? k1 = true *)
                     apply Nat.ltb_lt. exact H_k2_lt.
Qed.

(**
   Pairs in composed trace are pairwise compatible.

   Any two pairs in compose_trace T1 T2 are compatible.
   This follows from the transitivity of compatible_pairs.
*)
Lemma compose_trace_pairwise_compatible :
  forall (A B C : list Char) (T1 : Trace A B) (T2 : Trace B C)
         (p1 p2 : nat * nat),
    is_valid_trace_aux T1 = true ->
    is_valid_trace_aux T2 = true ->
    In p1 (compose_trace T1 T2) ->
    In p2 (compose_trace T1 T2) ->
    compatible_pairs p1 p2 = true.
Proof.
  intros A B C T1 T2 p1 p2 H_valid1 H_valid2 H_in1 H_in2.
  (* Destruct pairs to get components *)
  destruct p1 as [i1 k1].
  destruct p2 as [i2 k2].
  (* Extract witnesses for (i1, k1) using In_compose_trace *)
  apply In_compose_trace in H_in1 as [j1 [H_in1_T1 H_in1_T2]].
  (* Extract witnesses for (i2, k2) using In_compose_trace *)
  apply In_compose_trace in H_in2 as [j2 [H_in2_T1 H_in2_T2]].
  (* Apply transitivity of compatible_pairs *)
  eapply compatible_pairs_compose.
  - exact H_valid1.
  - exact H_valid2.
  - exact H_in1_T1.
  - exact H_in2_T1.
  - exact H_in1_T2.
  - exact H_in2_T2.
Qed.

(** * Phase 3: Trace Composition Cost Infrastructure *)

(** ** Sub-Phase 3.1: Touched Position Lemmas *)

(**
   Touched positions in A are preserved in composition.

   Positions touched in A by the composed trace are a subset of
   positions touched in A by T1.
*)
(**
   Helper: If i is in touched_in_A, then there exists k such that (i,k) is in the trace.
*)
Lemma In_touched_in_A_exists_pair :
  forall (A B : list Char) (T : Trace A B) (i : nat),
    In i (touched_in_A A B T) ->
    exists k, In (i, k) T.
Proof.
  intros A B T i H_in.
  induction T as [| [i' k'] T' IH].
  - simpl in H_in. contradiction.
  - simpl in H_in.
    destruct H_in as [H_eq | H_in'].
    + subst i. exists k'. left. reflexivity.
    + apply IH in H_in' as [k H_in_pair].
      exists k. right. exact H_in_pair.
Qed.

Lemma touched_in_A_incl :
  forall (A B C : list Char) (T1 : Trace A B) (T2 : Trace B C),
    incl (touched_in_A A C (compose_trace T1 T2)) (touched_in_A A B T1).
Proof.
  intros A B C T1 T2.
  unfold incl.
  intros i H_in.
  (* i is in touched_in_A of composed trace, so ∃k. (i,k) ∈ compose_trace T1 T2 *)
  apply In_touched_in_A_exists_pair in H_in as [k H_in_comp].
  (* By In_compose_trace, ∃j. (i,j)∈T1 ∧ (j,k)∈T2 *)
  apply In_compose_trace in H_in_comp as [j [H_in_T1 H_in_T2]].
  (* Now show i ∈ touched_in_A A B T1 *)
  clear H_in_T2 k.
  induction T1 as [| [i1 j1] T1' IH_T1].
  - simpl in H_in_T1. contradiction.
  - simpl in H_in_T1.
    destruct H_in_T1 as [H_eq_pair | H_in_T1'].
    + injection H_eq_pair as H_i H_j. subst i1.
      simpl. left. reflexivity.
    + simpl. right. apply IH_T1. exact H_in_T1'.
Qed.

(**
   Touched positions in B are preserved in composition.

   Positions touched in C by the composed trace are a subset of
   positions touched in C by T2.
*)
(**
   Helper: If k is in touched_in_B, then there exists i such that (i,k) is in the trace.
*)
Lemma In_touched_in_B_exists_pair :
  forall (A B : list Char) (T : Trace A B) (k : nat),
    In k (touched_in_B A B T) ->
    exists i, In (i, k) T.
Proof.
  intros A B T k H_in.
  induction T as [| [i' k'] T' IH].
  - simpl in H_in. contradiction.
  - simpl in H_in.
    destruct H_in as [H_eq | H_in'].
    + subst k. exists i'. left. reflexivity.
    + apply IH in H_in' as [i H_in_pair].
      exists i. right. exact H_in_pair.
Qed.

Lemma touched_in_B_incl :
  forall (A B C : list Char) (T1 : Trace A B) (T2 : Trace B C),
    incl (touched_in_B A C (compose_trace T1 T2)) (touched_in_B B C T2).
Proof.
  intros A B C T1 T2.
  unfold incl.
  intros k H_in.
  (* k is in touched_in_B of composed trace, so ∃i. (i,k) ∈ compose_trace T1 T2 *)
  apply In_touched_in_B_exists_pair in H_in as [i H_in_comp].
  (* By In_compose_trace, ∃j. (i,j)∈T1 ∧ (j,k)∈T2 *)
  apply In_compose_trace in H_in_comp as [j [H_in_T1 H_in_T2]].
  (* Now show k ∈ touched_in_B B C T2 *)
  clear H_in_T1 i.
  induction T2 as [| [j2 k2] T2' IH_T2].
  - simpl in H_in_T2. contradiction.
  - simpl in H_in_T2.
    destruct H_in_T2 as [H_eq_pair | H_in_T2'].
    + injection H_eq_pair as H_j H_k. subst k2.
      simpl. left. reflexivity.
    + simpl. right. apply IH_T2. exact H_in_T2'.
Qed.

(**
   Substitution cost is bounded by 1.
*)
Lemma subst_cost_bound :
  forall c1 c2 : Char, subst_cost c1 c2 <= 1.
Proof.
  intros c1 c2.
  unfold subst_cost.
  destruct (char_eq c1 c2); lia.
Qed.

(**
   If l1 is included in l2, then length l1 ≤ length l2.

   Note: This is a general list property, may already exist in stdlib.
*)
Lemma incl_length :
  forall {A : Type} (l1 l2 : list A),
    incl l1 l2 ->
    NoDup l2 ->
    length l1 <= length l2.
Proof.
  intros A l1 l2 H_incl H_nodup.
  (* This requires counting elements, which is non-trivial without NoDup on l1 *)
  (* For now, we'll use a weaker approach that works even with duplicates in l1 *)
  induction l1 as [| a l1' IH].
  - (* Base: l1 = [] *)
    simpl. lia.
  - (* Inductive: l1 = a :: l1' *)
    simpl.
    (* We need: 1 + length l1' ≤ length l2 *)
    (* By H_incl, a ∈ l2, so length l2 ≥ 1 *)
    (* Also incl l1' l2, so by IH, length l1' ≤ length l2 *)
    (* But this doesn't directly give us what we need without NoDup on l1 *)
    (* Let's admit this for now and come back if needed *)
    admit.
Admitted.

(** ** Sub-Phase 3.2: Change Cost Infrastructure *)

(**
   Substitution cost satisfies weak triangle inequality.

   The cost of substituting a for c is at most the cost of substituting
   a for b plus the cost of substituting b for c.
*)
Lemma subst_cost_triangle :
  forall (a b c : Char),
    subst_cost a c <= subst_cost a b + subst_cost b c.
Proof.
  intros a b c.
  unfold subst_cost.
  destruct (char_eq a b) eqn:Eab;
  destruct (char_eq b c) eqn:Ebc;
  destruct (char_eq a c) eqn:Eac; simpl; try lia;
  (* Three impossible cases remain - all involve transitivity contradictions *)
  repeat match goal with
  | H1: char_eq ?x ?y = true, H2: char_eq ?y ?z = true |- _ =>
      apply char_eq_correct in H1; apply char_eq_correct in H2; subst
  end;
  match goal with
  | H: char_eq ?x ?x = false |- _ =>
      assert (Hrefl: char_eq x x = true) by (apply char_eq_correct; reflexivity);
      rewrite Hrefl in H; discriminate
  end.
Qed.

(**
   Length of touched positions is bounded by trace length.

   Each pair in the trace contributes one position to touched_in_A.
*)
Lemma touched_length_bound_A :
  forall (A B : list Char) (T : Trace A B),
    length (touched_in_A A B T) <= length T.
Proof.
  intros A B T.
  induction T as [| [i j] T' IH].
  - (* Base: T = [] *)
    simpl. lia.
  - (* Inductive: T = (i,j) :: T' *)
    simpl.
    lia.
Qed.

(**
   Length of touched positions in B is bounded by trace length.

   Each pair in the trace contributes one position to touched_in_B.
*)
Lemma touched_length_bound_B :
  forall (A B : list Char) (T : Trace A B),
    length (touched_in_B A B T) <= length T.
Proof.
  intros A B T.
  induction T as [| [i j] T' IH].
  - (* Base: T = [] *)
    simpl. lia.
  - (* Inductive: T = (i,j) :: T' *)
    simpl.
    lia.
Qed.

(**
   Trace Composition Preserves Validity

   If T1 is a valid trace from A to B and T2 is a valid trace from B to C,
   then their composition T1∘T2 is a valid trace from A to C.

   A valid trace must satisfy:
   1. All pairs have valid positions (1 ≤ i ≤ |A|, 1 ≤ k ≤ |C|)
   2. Pairs are compatible (no crossing lines, at most one match per position)

   Proof strategy:
   - Show composed pairs (i,k) have valid positions by transitivity
   - Show order preservation: if (i₁,j₁) and (j₁,k₁) ∈ T1∘T2, and (i₂,j₂) and (j₂,k₂) ∈ T1∘T2,
     then i₁ < i₂ ⟺ j₁ < j₂ and j₁ < j₂ ⟺ k₁ < k₂, thus i₁ < i₂ ⟺ k₁ < k₂
   - Show each position touched at most once follows from same property in T1 and T2
*)
Lemma compose_trace_preserves_validity :
  forall (A B C : list Char) (T1 : Trace A B) (T2 : Trace B C),
    is_valid_trace A B T1 = true ->
    is_valid_trace B C T2 = true ->
    is_valid_trace A C (compose_trace T1 T2) = true.
Proof.
  intros A B C T1 T2 H_valid1 H_valid2.
  unfold is_valid_trace in *.
  rewrite andb_true_iff in *.
  destruct H_valid1 as [H_bounds1 H_compat1].
  destruct H_valid2 as [H_bounds2 H_compat2].
  split.

  - (* Part 1: All pairs in composed trace have valid bounds *)
    apply forallb_forall.
    intros [i k] H_in.
    rewrite In_compose_trace in H_in.
    destruct H_in as [j [H_in1 H_in2]].
    (* Use valid_pair_compose with witnesses *)
    rewrite forallb_forall in H_bounds1.
    rewrite forallb_forall in H_bounds2.
    apply valid_pair_compose with (lenB := length B) (j := j).
    + apply H_bounds1. exact H_in1.
    + apply H_bounds2. exact H_in2.

  - (* Part 2: All pairs in composed trace are pairwise compatible *)
    (* Build is_valid_trace_aux from pairwise compatibility *)
    apply is_valid_trace_aux_from_pairwise.
    intros p1 p2 H_in1 H_in2.
    (* Use compose_trace_pairwise_compatible with the helper lemmas *)
    eapply compose_trace_pairwise_compatible.
    + exact H_compat1.
    + exact H_compat2.
    + exact H_in1.
    + exact H_in2.
Qed.

(** ** Sub-Phase 3.3: Change Cost Bound *)

(**
   Change Cost Composition Bound

   The change cost of a composed trace is bounded by the sum of change costs
   from the individual traces.

   ADMITTED - Requires fold_left infrastructure (deferred to Phase 4)

   Proof Strategy:
   For each pair (i,k) in compose_trace T1 T2:
   1. Use In_compose_trace to extract witness j such that (i,j)∈T1 and (j,k)∈T2
   2. Apply subst_cost_triangle:
      subst_cost(A[i-1], C[k-1]) ≤ subst_cost(A[i-1], B[j-1]) + subst_cost(B[j-1], C[k-1])
   3. Sum over all pairs in the composition using fold_left monotonicity

   Required Infrastructure (Phase 4):
   - fold_left_add_monotone: If f p ≤ g p pointwise, then fold_left adds preserve ≤
   - pair_cost_witness: For each pair in composition, construct witness pair in T1×T2
   - sum_bound_from_pointwise: Summation of fold_left preserves pointwise inequalities

   Key Challenge:
   The composition may have multiple pairs sharing the same witness in T1 or T2,
   so we need careful handling of multiplicity in the sum.

   Alternative Approaches:
   - Direct induction on structure of compose_trace (awkward due to fold_left definition)
   - Build general theory of fold_left summation with witness functions
   - Use list inclusion properties to bound sums (current planned approach)

   Estimated Complexity: ~60-80 lines
   Estimated Time: ~3-4 hours

   Note: This lemma is the main technical obstacle in Phase 3. Everything else
   (including the triangle inequality proof) works once this is proven.
*)
Lemma change_cost_compose_bound :
  forall (A B C : list Char) (T1 : Trace A B) (T2 : Trace B C),
    fold_left (fun acc p =>
      let '(i, k) := p in
      acc + subst_cost (nth (i-1) A default_char) (nth (k-1) C default_char)
    ) (compose_trace T1 T2) 0
    <=
    fold_left (fun acc p =>
      let '(i, j) := p in
      acc + subst_cost (nth (i-1) A default_char) (nth (j-1) B default_char)
    ) T1 0 +
    fold_left (fun acc p =>
      let '(j, k) := p in
      acc + subst_cost (nth (j-1) B default_char) (nth (k-1) C default_char)
    ) T2 0.
Proof.
  (* TODO Phase 4: Requires fold_left summation infrastructure *)
  admit.
Admitted.

(** ** Sub-Phase 3.4: Main Theorem *)

(**
   Lemma 1 (Wagner-Fischer, 1974, page 3):
   Trace Composition Cost Bound

   The cost of a composed trace is at most the sum of the individual trace costs.
   This is the key lemma enabling the triangle inequality proof.

   Intuition:
   - If position i in A is matched to j in B (by T1), and j in B is matched to k in C (by T2),
     then in the composed trace T1∘T2, position i in A is matched directly to k in C
   - The change cost in the composition is at most the sum of change costs from both traces
   - Positions touched in intermediate string B but not matched in composition become
     deletions from A and insertions to C, counted in both original costs

   This proof requires careful accounting of:
   1. Which positions are touched in each string
   2. How matched pairs contribute to change costs
   3. How unmatched positions contribute to insertion/deletion costs
*)
Lemma trace_composition_cost_bound :
  forall (A B C : list Char) (T1 : Trace A B) (T2 : Trace B C),
    trace_cost A C (compose_trace T1 T2) <= trace_cost A B T1 + trace_cost B C T2.
Proof.
  intros A B C T1 T2.
  unfold trace_cost.

  (* Introduce convenient notation for the three cost components of each trace *)
  set (comp := compose_trace T1 T2).
  set (cc_comp := fold_left (fun acc p =>
    let '(i, k) := p in
    acc + subst_cost (nth (i-1) A default_char) (nth (k-1) C default_char)
  ) comp 0).
  set (dc_comp := length A - length (touched_in_A A C comp)).
  set (ic_comp := length C - length (touched_in_B A C comp)).

  set (cc1 := fold_left (fun acc p =>
    let '(i, j) := p in
    acc + subst_cost (nth (i-1) A default_char) (nth (j-1) B default_char)
  ) T1 0).
  set (dc1 := length A - length (touched_in_A A B T1)).
  set (ic1 := length B - length (touched_in_B A B T1)).

  set (cc2 := fold_left (fun acc p =>
    let '(j, k) := p in
    acc + subst_cost (nth (j-1) B default_char) (nth (k-1) C default_char)
  ) T2 0).
  set (dc2 := length B - length (touched_in_A B C T2)).
  set (ic2 := length C - length (touched_in_B B C T2)).

  (* Goal: cc_comp + dc_comp + ic_comp <= (cc1 + dc1 + ic1) + (cc2 + dc2 + ic2) *)

  (* Part 1: Bound change costs using triangle inequality *)
  assert (H_cc: cc_comp <= cc1 + cc2).
  { unfold cc_comp, cc1, cc2, comp.
    apply change_cost_compose_bound.
  }

  (* Part 2: Bound delete + insert costs using the 2|B| slack *)
  (* This is where the 2|B| term provides slack to make the inequality work *)
  (* For Phase 3, we observe that this bound holds but defer the full arithmetic proof to Phase 4 *)
  assert (H_di: dc_comp + ic_comp <= dc1 + ic1 + dc2 + ic2).
  { unfold dc_comp, ic_comp, dc1, ic1, dc2, ic2, comp.
    (* TODO Phase 4: Rigorous proof of delete/insert cost bound using 2|B| slack *)
    admit.
  }

  (* Combine the two bounds *)
  lia.
Admitted.

(**
   Theorem 1 (Wagner-Fischer, 1974, page 4):
   Distance-Trace Equivalence

   The recursive Levenshtein distance equals the minimum cost over all valid traces.

   This theorem bridges the recursive definition (which we've been working with)
   and the trace abstraction (which makes the triangle inequality trivial).

   Proof outline:
   1. Show that every valid trace corresponds to an edit sequence with the same cost
   2. Show that the optimal edit sequence corresponds to a trace with minimum cost
   3. Conclude equality

   This requires:
   - Proving the recursive definition computes minimum cost edit sequences
   - Proving trace cost accurately reflects edit operation costs
   - Showing the correspondence is bijective for optimal solutions
*)
Theorem distance_equals_min_trace_cost :
  forall (A B : list Char),
    exists (T_opt : Trace A B),
      is_valid_trace A B T_opt = true /\
      trace_cost A B T_opt = lev_distance A B /\
      (forall T : Trace A B, is_valid_trace A B T = true ->
        trace_cost A B T_opt <= trace_cost A B T).
Proof.
  intros A B.
  (* This theorem requires:
     1. Constructing an optimal trace from the recursive distance computation
     2. Proving this trace has cost equal to lev_distance
     3. Proving it's minimal among all valid traces

     Strategy:
     - Use the DP matrix to extract an optimal trace (backtracking)
     - Prove the trace is valid
     - Prove its cost equals the distance
     - Prove optimality by showing any cheaper trace would contradict the DP recurrence

     This is a substantial proof that requires formalizing:
     - Trace extraction from DP matrix
     - Trace validity preservation
     - Cost equivalence

     For now, we admit this and use it to prove the triangle inequality,
     then return to complete this proof.
  *)
  admit.
Admitted.

(** Theorem: Triangle inequality - distance satisfies metric property *)
(**
   Proof Strategy (Wagner-Fischer 1974):

   Instead of complex induction on intermediate strings with nested min3 expressions,
   we use the trace abstraction and prove via trace composition.

   Key insights:
   1. Theorem 1: d(A, B) = min{cost(T) | T: A→B is valid}
   2. Lemma 1: cost(T₁ ∘ T₂) ≤ cost(T₁) + cost(T₂)

   From this, the triangle inequality follows immediately:
     d(A, C) = min{cost(T) | T: A→C}                    [by Theorem 1]
            ≤ cost(T₁ ∘ T₂)                              [for optimal T₁: A→B, T₂: B→C]
            ≤ cost(T₁) + cost(T₂)                        [by Lemma 1]
            = d(A, B) + d(B, C)                          [by Theorem 1]
*)
Theorem lev_distance_triangle_inequality :
  forall (s1 s2 s3 : list Char),
    lev_distance s1 s3 <= lev_distance s1 s2 + lev_distance s2 s3.
Proof.
  intros s1 s2 s3.

  (* By Theorem 1, there exist optimal traces T1: s1→s2 and T2: s2→s3 *)
  destruct (distance_equals_min_trace_cost s1 s2) as [T1 [H_valid1 [H_cost1 H_opt1]]].
  destruct (distance_equals_min_trace_cost s2 s3) as [T2 [H_valid2 [H_cost2 H_opt2]]].

  (* Compose the traces: T_comp = T1 ∘ T2 : s1→s3 *)
  set (T_comp := compose_trace T1 T2).

  (* By Theorem 1, there exists an optimal trace for s1→s3 *)
  destruct (distance_equals_min_trace_cost s1 s3) as [T_opt [H_valid_opt [H_cost_opt H_opt]]].

  (* Now we show: d(s1,s3) ≤ d(s1,s2) + d(s2,s3) *)
  rewrite <- H_cost_opt.           (* d(s1,s3) = cost(T_opt) *)
  rewrite <- H_cost1.              (* d(s1,s2) = cost(T1) *)
  rewrite <- H_cost2.              (* d(s2,s3) = cost(T2) *)

  (* Need to prove: cost(T_opt) ≤ cost(T1) + cost(T2) *)

  (* Prove that T_comp is valid using compose_trace_preserves_validity *)
  assert (H_comp_valid: is_valid_trace s1 s3 T_comp = true).
  {
    unfold T_comp.
    apply compose_trace_preserves_validity.
    - exact H_valid1.
    - exact H_valid2.
  }

  (* By optimality of T_opt, we have cost(T_opt) ≤ cost(T_comp) *)
  assert (H_bound: trace_cost s1 s3 T_opt <= trace_cost s1 s3 T_comp).
  {
    apply H_opt.
    exact H_comp_valid.
  }

  (* By Lemma 1, we have cost(T_comp) ≤ cost(T1) + cost(T2) *)
  assert (H_lemma1: trace_cost s1 s3 T_comp <= trace_cost s1 s2 T1 + trace_cost s2 s3 T2).
  {
    unfold T_comp.
    apply trace_composition_cost_bound.
  }

  (* Combining the bounds: cost(T_opt) ≤ cost(T_comp) ≤ cost(T1) + cost(T2) *)
  lia.
Qed.

(*
(* ========================================================================== *)
(* ORIGINAL PARTIAL PROOF OF TRIANGLE INEQUALITY (saved for reference)       *)
(* This proof is incomplete and commented out. Left here for future reference *)
(* when completing the proof using well-founded induction.                    *)
(* ========================================================================== *)
(*
Proof.
  (* Key insight: Any edit sequence s1→s2→s3 is a valid (possibly suboptimal)
     edit sequence s1→s3. Since lev_distance computes the MINIMUM length
     sequence, the direct path s1→s3 cannot be longer than the concatenated
     path s1→s2→s3.

     Proof strategy: Induction on s2 (the intermediate string).
     This avoids needing to formalize full edit sequences while still
     capturing the composition property.

     Base case: s2 = [] means we go s1→[]→s3, which costs |s1| + |s3|.
                The direct path d(s1,s3) ≤ max(|s1|,|s3|) < |s1|+|s3|.

     Inductive step: s2 = c::s2', assume triangle inequality holds for s2',
                     show it holds for c::s2'. *)

  intros s1 s2 s3.

  (* Induction on s2 *)
  generalize dependent s3.
  generalize dependent s1.
  induction s2 as [| c2 s2' IHs2].

  - (* Base case: s2 = [] *)
    intros s1 s3.
    rewrite lev_distance_empty_left.
    rewrite lev_distance_empty_right.
    (* Need: d(s1, s3) ≤ |s1| + |s3| *)
    assert (H_upper: lev_distance s1 s3 <= Nat.max (length s1) (length s3)).
    { apply lev_distance_upper_bound. }
    lia.

  - (* Inductive case: s2 = c2 :: s2' *)
    intros s1 s3.
    (* IHs2: forall s1 s3, d(s1,s3) ≤ d(s1,s2') + d(s2',s3) *)

    (* Case analysis on s1 and s3 *)
    destruct s1 as [| c1 s1'].

    + (* s1 = [] *)
      (* d([],s3) ≤ d([],c2::s2') + d(c2::s2',s3) *)
      rewrite lev_distance_empty_left.
      (* |s3| ≤ d([],c2::s2') + d(c2::s2',s3) *)
      rewrite lev_distance_empty_left.
      (* |s3| ≤ |c2::s2'| + d(c2::s2',s3) *)
      (* Since d(c2::s2',s3) ≥ 0, this is true if |s3| ≤ |c2::s2'| + |s3| - |s3| *)
      (* Actually, we need |s3| ≤ S|s2'| + d(c2::s2',s3) *)
      (* Use: d(c2::s2',s3) ≥ abs(|c2::s2'| - |s3|) would give us this, but we don't have that *)
      (* Instead: |s3| ≤ S|s2'| + d(c2::s2',s3) is equivalent to needing d(c2::s2',s3) ≥ |s3| - S|s2'| *)
      (*This is just a fact about distance - we always need at least |difference in lengths| *)

      (* More direct: use that a ≤ b + c  if we know something about a, b, c *)
      simpl length.
      (* |s3| ≤ S|s2'| + d(c2::s2',s3) *)
      (* If |s3| ≤ S|s2'|, then this is trivial. Otherwise, d must compensate. *)
      (* Since we don't have the length-difference lemma proven, let's use the fact that
         the sum is at least max, and we know d(c2::s2',s3) is optimal. *)
      assert (H_case: length s3 <= S (length s2') \/ S (length s2') < length s3) by lia.
      destruct H_case as [H_s3_small | H_s3_large].
      * (* |s3| ≤ S|s2'| *)
        (* Then |s3| ≤ S|s2'| ≤ S|s2'| + d(c2::s2',s3) since d ≥ 0 *)
        transitivity (S (length s2')).
        { exact H_s3_small. }
        { apply Nat.le_add_r. }
      * (* S|s2'| < |s3| *)
        (* Then |s3| - S|s2'| > 0, and we need d(c2::s2',s3) ≥ |s3| - S|s2'| *)
        (* This is the length-difference lower bound, which we haven't proven *)
        (* For now, use upper bound theorem *)
        assert (H_upper: lev_distance (c2 :: s2') s3 <= Nat.max (S (length s2')) (length s3)).
        { apply lev_distance_upper_bound. }
        assert (H_max: Nat.max (S (length s2')) (length s3) = length s3).
        { apply Nat.max_r. lia. }
        rewrite H_max in H_upper.
        lia.

    + (* s1 = c1 :: s1' *)
      destruct s3 as [| c3 s3'].

      * (* s3 = [] *)
        rewrite lev_distance_empty_right.
        rewrite lev_distance_empty_right.
        (* Need: |c1::s1'| ≤ d(c1::s1', c2::s2') + |c2::s2'| *)
        assert (H_nonneg: 0 <= lev_distance (c1 :: s1') (c2 :: s2')).
        { lia. }
        lia.

      * (* s3 = c3 :: s3' *)
        (* All strings non-empty, use recursive definition *)
        rewrite lev_distance_cons.
        rewrite (lev_distance_cons c1 c2 s1' s2').
        rewrite (lev_distance_cons c2 c3 s2' s3').

        (* Now we have:
           min3 (d(s1',c3::s3')+1) (d(c1::s1',s3')+1) (d(s1',s3')+subst(c1,c3))
           ≤ min3 (d(s1',c2::s2')+1) (d(c1::s1',s2')+1) (d(s1',s2')+subst(c1,c2))
             + min3 (d(s2',c3::s3')+1) (d(c2::s2',s3')+1) (d(s2',s3')+subst(c2,c3))

           We'll show each branch of the LHS min3 is bounded by the RHS sum. *)

        (* Key insight: We can bound each case using IH on s2' *)
        assert (IH1: lev_distance s1' s3' <= lev_distance s1' s2' + lev_distance s2' s3').
        { apply IHs2. }
        assert (IH2: lev_distance s1' (c3 :: s3') <= lev_distance s1' s2' + lev_distance s2' (c3 :: s3')).
        { apply IHs2. }
        assert (IH3: lev_distance (c1 :: s1') s3' <= lev_distance (c1 :: s1') s2' + lev_distance s2' s3').
        { apply IHs2. }
        assert (IH4: lev_distance s1' (c3 :: s3') <= lev_distance s1' (c2 :: s2') + lev_distance (c2 :: s2') (c3 :: s3')).
        { apply IHs2. }
        assert (IH5: lev_distance (c1 :: s1') s3' <= lev_distance (c1 :: s1') (c2 :: s2') + lev_distance (c2 :: s2') s3').
        { apply IHs2. }

        (* Subst costs are bounded by 1 *)
        assert (H_subst_c1_c2: subst_cost c1 c2 <= 1).
        { unfold subst_cost. destruct (char_eq c1 c2); lia. }
        assert (H_subst_c2_c3: subst_cost c2 c3 <= 1).
        { unfold subst_cost. destruct (char_eq c2 c3); lia. }
        assert (H_subst_c1_c3: subst_cost c1 c3 <= 1).
        { unfold subst_cost. destruct (char_eq c1 c3); lia. }

        (* Use properties of min3 and the induction hypotheses *)
        unfold min3.

        (* The proof: min of LHS ≤ sum of RHS
           We show LHS ≤ RHS by showing each component of LHS min
           can be bounded by components of RHS. *)

        (* This requires careful arithmetic reasoning *)
        lia.
Qed.
*)
*)

(** * Main Correctness Theorem *)

(** This theorem states that IF a matrix is filled according to the
    Wagner-Fischer recurrence relation, THEN the value at position (i,j)
    equals the recursive Levenshtein distance between the first i and j
    characters of the input strings.

    The full proof of this theorem requires:
    1. Proper formalization of matrix filling (iterative loops)
    2. Strong induction on i + j
    3. Careful bookkeeping of matrix invariants

    This is substantial work and is admitted for now. *)
Theorem dp_matrix_correctness :
  forall (s1 s2 : list Char) (m : Matrix nat) (i j : nat),
    (* Preconditions: matrix properly initialized and filled *)
    i <= length s1 ->
    j <= length s2 ->
    (* If matrix follows Wagner-Fischer recurrence... *)
    (forall i' j',
      i' > 0 -> j' > 0 -> i' <= i -> j' <= j ->
      get_cell m i' j' = min3
        (get_cell m (i'-1) j' + 1)
        (get_cell m i' (j'-1) + 1)
        (get_cell m (i'-1) (j'-1) + subst_cost (nth (i'-1) s1 " "%char) (nth (j'-1) s2 " "%char))) ->
    (* Base cases *)
    (forall k, k <= i -> get_cell m k 0 = k) ->
    (forall k, k <= j -> get_cell m 0 k = k) ->
    (* Then matrix cell equals recursive distance *)
    get_cell m i j = lev_distance (firstn i s1) (firstn j s2).
Proof.
  (* This proof proceeds by strong induction on i + j, carefully applying
     the recurrence relation and induction hypothesis.

     It's the core correctness proof for the DP algorithm and requires
     significant detail. Admitted for now. *)
Admitted.

(** Helper lemma: firstn of full length is identity *)
Lemma firstn_all :
  forall {A : Type} (l : list A),
    firstn (length l) l = l.
Proof.
  intros A l.
  induction l as [| x xs IH].
  - simpl. reflexivity.
  - simpl. rewrite IH. reflexivity.
Qed.

(** * Corollary: Full Algorithm Correctness *)

(** When the matrix is fully computed for strings s1 and s2, the bottom-right
    cell contains the correct Levenshtein distance. *)
Corollary levenshtein_distance_correctness :
  forall (s1 s2 : list Char) (m : Matrix nat),
    (* If matrix is properly filled... *)
    (forall i j,
      i > 0 -> j > 0 -> i <= length s1 -> j <= length s2 ->
      get_cell m i j = min3
        (get_cell m (i-1) j + 1)
        (get_cell m i (j-1) + 1)
        (get_cell m (i-1) (j-1) + subst_cost (nth (i-1) s1 " "%char) (nth (j-1) s2 " "%char))) ->
    (forall k, k <= length s1 -> get_cell m k 0 = k) ->
    (forall k, k <= length s2 -> get_cell m 0 k = k) ->
    (* Then the final cell equals the recursive distance *)
    get_cell m (length s1) (length s2) = lev_distance s1 s2.
Proof.
  intros s1 s2 m H_recurrence H_row0 H_col0.

  (* Apply dp_matrix_correctness with i = length s1, j = length s2 *)
  assert (H_correct := dp_matrix_correctness s1 s2 m (length s1) (length s2)).

  (* Simplify H_correct using firstn_all *)
  rewrite !firstn_all in H_correct.

  apply H_correct.
  - lia.
  - lia.
  - intros i' j' H_i'_pos H_j'_pos H_i'_le H_j'_le.
    apply H_recurrence; lia.
  - exact H_row0.
  - exact H_col0.
Qed.

(** * Summary

    This module establishes the correctness of the Levenshtein distance algorithm:

    1. **Identity**: lev_distance s s = 0 ✓ PROVEN
    2. **Symmetry**: lev_distance s1 s2 = lev_distance s2 s1 (admitted)
    3. **Triangle inequality**: lev_distance s1 s3 ≤ lev_distance s1 s2 + lev_distance s2 s3 (admitted)
    4. **Upper bound**: lev_distance s1 s2 ≤ max(|s1|, |s2|) (admitted)
    5. **DP correctness**: Matrix algorithm equals recursive definition (admitted)

    The admitted proofs are standard results in edit distance theory and can be
    completed following well-established proof techniques. The infrastructure
    (definitions, basic lemmas, proof structure) is in place for completing them.
*)
